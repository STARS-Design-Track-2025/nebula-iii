module team_05 (ACK_I,
    CYC_O,
    STB_O,
    WE_O,
    clk,
    en,
    nrst,
    vccd1,
    vssd1,
    ADR_O,
    DAT_I,
    DAT_O,
    SEL_O,
    gpio_in,
    gpio_oeb,
    gpio_out);
 input ACK_I;
 output CYC_O;
 output STB_O;
 output WE_O;
 input clk;
 input en;
 input nrst;
 input vccd1;
 input vssd1;
 output [31:0] ADR_O;
 input [31:0] DAT_I;
 output [31:0] DAT_O;
 output [3:0] SEL_O;
 input [33:0] gpio_in;
 output [33:0] gpio_oeb;
 output [33:0] gpio_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire clknet_leaf_0_clk;
 wire \top.CB_read_complete ;
 wire \top.CB_write_complete ;
 wire \top.FLV_done ;
 wire \top.HT_fin_reg ;
 wire \top.TRN_char_index[0] ;
 wire \top.TRN_char_index[1] ;
 wire \top.TRN_char_index[2] ;
 wire \top.TRN_char_index[3] ;
 wire \top.TRN_char_index[4] ;
 wire \top.TRN_char_index[5] ;
 wire \top.TRN_char_index[6] ;
 wire \top.TRN_sram_complete ;
 wire \top.WB.CPU_DAT_O[0] ;
 wire \top.WB.CPU_DAT_O[10] ;
 wire \top.WB.CPU_DAT_O[11] ;
 wire \top.WB.CPU_DAT_O[12] ;
 wire \top.WB.CPU_DAT_O[13] ;
 wire \top.WB.CPU_DAT_O[14] ;
 wire \top.WB.CPU_DAT_O[15] ;
 wire \top.WB.CPU_DAT_O[16] ;
 wire \top.WB.CPU_DAT_O[17] ;
 wire \top.WB.CPU_DAT_O[18] ;
 wire \top.WB.CPU_DAT_O[19] ;
 wire \top.WB.CPU_DAT_O[1] ;
 wire \top.WB.CPU_DAT_O[20] ;
 wire \top.WB.CPU_DAT_O[21] ;
 wire \top.WB.CPU_DAT_O[22] ;
 wire \top.WB.CPU_DAT_O[23] ;
 wire \top.WB.CPU_DAT_O[24] ;
 wire \top.WB.CPU_DAT_O[25] ;
 wire \top.WB.CPU_DAT_O[26] ;
 wire \top.WB.CPU_DAT_O[27] ;
 wire \top.WB.CPU_DAT_O[28] ;
 wire \top.WB.CPU_DAT_O[29] ;
 wire \top.WB.CPU_DAT_O[2] ;
 wire \top.WB.CPU_DAT_O[30] ;
 wire \top.WB.CPU_DAT_O[31] ;
 wire \top.WB.CPU_DAT_O[3] ;
 wire \top.WB.CPU_DAT_O[4] ;
 wire \top.WB.CPU_DAT_O[5] ;
 wire \top.WB.CPU_DAT_O[6] ;
 wire \top.WB.CPU_DAT_O[7] ;
 wire \top.WB.CPU_DAT_O[8] ;
 wire \top.WB.CPU_DAT_O[9] ;
 wire \top.WB.curr_state[0] ;
 wire \top.WB.curr_state[1] ;
 wire \top.WB.curr_state[2] ;
 wire \top.WB.prev_BUSY_O ;
 wire \top.WorR ;
 wire \top.cb_syn.cb_enable ;
 wire \top.cb_syn.cb_length[0] ;
 wire \top.cb_syn.cb_length[1] ;
 wire \top.cb_syn.cb_length[2] ;
 wire \top.cb_syn.cb_length[3] ;
 wire \top.cb_syn.cb_length[4] ;
 wire \top.cb_syn.cb_length[5] ;
 wire \top.cb_syn.cb_length[6] ;
 wire \top.cb_syn.char_found ;
 wire \top.cb_syn.char_index[0] ;
 wire \top.cb_syn.char_index[1] ;
 wire \top.cb_syn.char_index[2] ;
 wire \top.cb_syn.char_index[3] ;
 wire \top.cb_syn.char_index[4] ;
 wire \top.cb_syn.char_index[5] ;
 wire \top.cb_syn.char_index[6] ;
 wire \top.cb_syn.char_index[7] ;
 wire \top.cb_syn.char_path[0] ;
 wire \top.cb_syn.char_path[100] ;
 wire \top.cb_syn.char_path[101] ;
 wire \top.cb_syn.char_path[102] ;
 wire \top.cb_syn.char_path[103] ;
 wire \top.cb_syn.char_path[104] ;
 wire \top.cb_syn.char_path[105] ;
 wire \top.cb_syn.char_path[106] ;
 wire \top.cb_syn.char_path[107] ;
 wire \top.cb_syn.char_path[108] ;
 wire \top.cb_syn.char_path[109] ;
 wire \top.cb_syn.char_path[10] ;
 wire \top.cb_syn.char_path[110] ;
 wire \top.cb_syn.char_path[111] ;
 wire \top.cb_syn.char_path[112] ;
 wire \top.cb_syn.char_path[113] ;
 wire \top.cb_syn.char_path[114] ;
 wire \top.cb_syn.char_path[115] ;
 wire \top.cb_syn.char_path[116] ;
 wire \top.cb_syn.char_path[117] ;
 wire \top.cb_syn.char_path[118] ;
 wire \top.cb_syn.char_path[119] ;
 wire \top.cb_syn.char_path[11] ;
 wire \top.cb_syn.char_path[120] ;
 wire \top.cb_syn.char_path[121] ;
 wire \top.cb_syn.char_path[122] ;
 wire \top.cb_syn.char_path[123] ;
 wire \top.cb_syn.char_path[124] ;
 wire \top.cb_syn.char_path[125] ;
 wire \top.cb_syn.char_path[126] ;
 wire \top.cb_syn.char_path[127] ;
 wire \top.cb_syn.char_path[12] ;
 wire \top.cb_syn.char_path[13] ;
 wire \top.cb_syn.char_path[14] ;
 wire \top.cb_syn.char_path[15] ;
 wire \top.cb_syn.char_path[16] ;
 wire \top.cb_syn.char_path[17] ;
 wire \top.cb_syn.char_path[18] ;
 wire \top.cb_syn.char_path[19] ;
 wire \top.cb_syn.char_path[1] ;
 wire \top.cb_syn.char_path[20] ;
 wire \top.cb_syn.char_path[21] ;
 wire \top.cb_syn.char_path[22] ;
 wire \top.cb_syn.char_path[23] ;
 wire \top.cb_syn.char_path[24] ;
 wire \top.cb_syn.char_path[25] ;
 wire \top.cb_syn.char_path[26] ;
 wire \top.cb_syn.char_path[27] ;
 wire \top.cb_syn.char_path[28] ;
 wire \top.cb_syn.char_path[29] ;
 wire \top.cb_syn.char_path[2] ;
 wire \top.cb_syn.char_path[30] ;
 wire \top.cb_syn.char_path[31] ;
 wire \top.cb_syn.char_path[32] ;
 wire \top.cb_syn.char_path[33] ;
 wire \top.cb_syn.char_path[34] ;
 wire \top.cb_syn.char_path[35] ;
 wire \top.cb_syn.char_path[36] ;
 wire \top.cb_syn.char_path[37] ;
 wire \top.cb_syn.char_path[38] ;
 wire \top.cb_syn.char_path[39] ;
 wire \top.cb_syn.char_path[3] ;
 wire \top.cb_syn.char_path[40] ;
 wire \top.cb_syn.char_path[41] ;
 wire \top.cb_syn.char_path[42] ;
 wire \top.cb_syn.char_path[43] ;
 wire \top.cb_syn.char_path[44] ;
 wire \top.cb_syn.char_path[45] ;
 wire \top.cb_syn.char_path[46] ;
 wire \top.cb_syn.char_path[47] ;
 wire \top.cb_syn.char_path[48] ;
 wire \top.cb_syn.char_path[49] ;
 wire \top.cb_syn.char_path[4] ;
 wire \top.cb_syn.char_path[50] ;
 wire \top.cb_syn.char_path[51] ;
 wire \top.cb_syn.char_path[52] ;
 wire \top.cb_syn.char_path[53] ;
 wire \top.cb_syn.char_path[54] ;
 wire \top.cb_syn.char_path[55] ;
 wire \top.cb_syn.char_path[56] ;
 wire \top.cb_syn.char_path[57] ;
 wire \top.cb_syn.char_path[58] ;
 wire \top.cb_syn.char_path[59] ;
 wire \top.cb_syn.char_path[5] ;
 wire \top.cb_syn.char_path[60] ;
 wire \top.cb_syn.char_path[61] ;
 wire \top.cb_syn.char_path[62] ;
 wire \top.cb_syn.char_path[63] ;
 wire \top.cb_syn.char_path[64] ;
 wire \top.cb_syn.char_path[65] ;
 wire \top.cb_syn.char_path[66] ;
 wire \top.cb_syn.char_path[67] ;
 wire \top.cb_syn.char_path[68] ;
 wire \top.cb_syn.char_path[69] ;
 wire \top.cb_syn.char_path[6] ;
 wire \top.cb_syn.char_path[70] ;
 wire \top.cb_syn.char_path[71] ;
 wire \top.cb_syn.char_path[72] ;
 wire \top.cb_syn.char_path[73] ;
 wire \top.cb_syn.char_path[74] ;
 wire \top.cb_syn.char_path[75] ;
 wire \top.cb_syn.char_path[76] ;
 wire \top.cb_syn.char_path[77] ;
 wire \top.cb_syn.char_path[78] ;
 wire \top.cb_syn.char_path[79] ;
 wire \top.cb_syn.char_path[7] ;
 wire \top.cb_syn.char_path[80] ;
 wire \top.cb_syn.char_path[81] ;
 wire \top.cb_syn.char_path[82] ;
 wire \top.cb_syn.char_path[83] ;
 wire \top.cb_syn.char_path[84] ;
 wire \top.cb_syn.char_path[85] ;
 wire \top.cb_syn.char_path[86] ;
 wire \top.cb_syn.char_path[87] ;
 wire \top.cb_syn.char_path[88] ;
 wire \top.cb_syn.char_path[89] ;
 wire \top.cb_syn.char_path[8] ;
 wire \top.cb_syn.char_path[90] ;
 wire \top.cb_syn.char_path[91] ;
 wire \top.cb_syn.char_path[92] ;
 wire \top.cb_syn.char_path[93] ;
 wire \top.cb_syn.char_path[94] ;
 wire \top.cb_syn.char_path[95] ;
 wire \top.cb_syn.char_path[96] ;
 wire \top.cb_syn.char_path[97] ;
 wire \top.cb_syn.char_path[98] ;
 wire \top.cb_syn.char_path[99] ;
 wire \top.cb_syn.char_path[9] ;
 wire \top.cb_syn.char_path_n[0] ;
 wire \top.cb_syn.char_path_n[100] ;
 wire \top.cb_syn.char_path_n[101] ;
 wire \top.cb_syn.char_path_n[102] ;
 wire \top.cb_syn.char_path_n[103] ;
 wire \top.cb_syn.char_path_n[104] ;
 wire \top.cb_syn.char_path_n[105] ;
 wire \top.cb_syn.char_path_n[106] ;
 wire \top.cb_syn.char_path_n[107] ;
 wire \top.cb_syn.char_path_n[108] ;
 wire \top.cb_syn.char_path_n[109] ;
 wire \top.cb_syn.char_path_n[10] ;
 wire \top.cb_syn.char_path_n[110] ;
 wire \top.cb_syn.char_path_n[111] ;
 wire \top.cb_syn.char_path_n[112] ;
 wire \top.cb_syn.char_path_n[113] ;
 wire \top.cb_syn.char_path_n[114] ;
 wire \top.cb_syn.char_path_n[115] ;
 wire \top.cb_syn.char_path_n[116] ;
 wire \top.cb_syn.char_path_n[117] ;
 wire \top.cb_syn.char_path_n[118] ;
 wire \top.cb_syn.char_path_n[119] ;
 wire \top.cb_syn.char_path_n[11] ;
 wire \top.cb_syn.char_path_n[120] ;
 wire \top.cb_syn.char_path_n[121] ;
 wire \top.cb_syn.char_path_n[122] ;
 wire \top.cb_syn.char_path_n[123] ;
 wire \top.cb_syn.char_path_n[124] ;
 wire \top.cb_syn.char_path_n[125] ;
 wire \top.cb_syn.char_path_n[126] ;
 wire \top.cb_syn.char_path_n[127] ;
 wire \top.cb_syn.char_path_n[12] ;
 wire \top.cb_syn.char_path_n[13] ;
 wire \top.cb_syn.char_path_n[14] ;
 wire \top.cb_syn.char_path_n[15] ;
 wire \top.cb_syn.char_path_n[16] ;
 wire \top.cb_syn.char_path_n[17] ;
 wire \top.cb_syn.char_path_n[18] ;
 wire \top.cb_syn.char_path_n[19] ;
 wire \top.cb_syn.char_path_n[1] ;
 wire \top.cb_syn.char_path_n[20] ;
 wire \top.cb_syn.char_path_n[21] ;
 wire \top.cb_syn.char_path_n[22] ;
 wire \top.cb_syn.char_path_n[23] ;
 wire \top.cb_syn.char_path_n[24] ;
 wire \top.cb_syn.char_path_n[25] ;
 wire \top.cb_syn.char_path_n[26] ;
 wire \top.cb_syn.char_path_n[27] ;
 wire \top.cb_syn.char_path_n[28] ;
 wire \top.cb_syn.char_path_n[29] ;
 wire \top.cb_syn.char_path_n[2] ;
 wire \top.cb_syn.char_path_n[30] ;
 wire \top.cb_syn.char_path_n[31] ;
 wire \top.cb_syn.char_path_n[32] ;
 wire \top.cb_syn.char_path_n[33] ;
 wire \top.cb_syn.char_path_n[34] ;
 wire \top.cb_syn.char_path_n[35] ;
 wire \top.cb_syn.char_path_n[36] ;
 wire \top.cb_syn.char_path_n[37] ;
 wire \top.cb_syn.char_path_n[38] ;
 wire \top.cb_syn.char_path_n[39] ;
 wire \top.cb_syn.char_path_n[3] ;
 wire \top.cb_syn.char_path_n[40] ;
 wire \top.cb_syn.char_path_n[41] ;
 wire \top.cb_syn.char_path_n[42] ;
 wire \top.cb_syn.char_path_n[43] ;
 wire \top.cb_syn.char_path_n[44] ;
 wire \top.cb_syn.char_path_n[45] ;
 wire \top.cb_syn.char_path_n[46] ;
 wire \top.cb_syn.char_path_n[47] ;
 wire \top.cb_syn.char_path_n[48] ;
 wire \top.cb_syn.char_path_n[49] ;
 wire \top.cb_syn.char_path_n[4] ;
 wire \top.cb_syn.char_path_n[50] ;
 wire \top.cb_syn.char_path_n[51] ;
 wire \top.cb_syn.char_path_n[52] ;
 wire \top.cb_syn.char_path_n[53] ;
 wire \top.cb_syn.char_path_n[54] ;
 wire \top.cb_syn.char_path_n[55] ;
 wire \top.cb_syn.char_path_n[56] ;
 wire \top.cb_syn.char_path_n[57] ;
 wire \top.cb_syn.char_path_n[58] ;
 wire \top.cb_syn.char_path_n[59] ;
 wire \top.cb_syn.char_path_n[5] ;
 wire \top.cb_syn.char_path_n[60] ;
 wire \top.cb_syn.char_path_n[61] ;
 wire \top.cb_syn.char_path_n[62] ;
 wire \top.cb_syn.char_path_n[63] ;
 wire \top.cb_syn.char_path_n[64] ;
 wire \top.cb_syn.char_path_n[65] ;
 wire \top.cb_syn.char_path_n[66] ;
 wire \top.cb_syn.char_path_n[67] ;
 wire \top.cb_syn.char_path_n[68] ;
 wire \top.cb_syn.char_path_n[69] ;
 wire \top.cb_syn.char_path_n[6] ;
 wire \top.cb_syn.char_path_n[70] ;
 wire \top.cb_syn.char_path_n[71] ;
 wire \top.cb_syn.char_path_n[72] ;
 wire \top.cb_syn.char_path_n[73] ;
 wire \top.cb_syn.char_path_n[74] ;
 wire \top.cb_syn.char_path_n[75] ;
 wire \top.cb_syn.char_path_n[76] ;
 wire \top.cb_syn.char_path_n[77] ;
 wire \top.cb_syn.char_path_n[78] ;
 wire \top.cb_syn.char_path_n[79] ;
 wire \top.cb_syn.char_path_n[7] ;
 wire \top.cb_syn.char_path_n[80] ;
 wire \top.cb_syn.char_path_n[81] ;
 wire \top.cb_syn.char_path_n[82] ;
 wire \top.cb_syn.char_path_n[83] ;
 wire \top.cb_syn.char_path_n[84] ;
 wire \top.cb_syn.char_path_n[85] ;
 wire \top.cb_syn.char_path_n[86] ;
 wire \top.cb_syn.char_path_n[87] ;
 wire \top.cb_syn.char_path_n[88] ;
 wire \top.cb_syn.char_path_n[89] ;
 wire \top.cb_syn.char_path_n[8] ;
 wire \top.cb_syn.char_path_n[90] ;
 wire \top.cb_syn.char_path_n[91] ;
 wire \top.cb_syn.char_path_n[92] ;
 wire \top.cb_syn.char_path_n[93] ;
 wire \top.cb_syn.char_path_n[94] ;
 wire \top.cb_syn.char_path_n[95] ;
 wire \top.cb_syn.char_path_n[96] ;
 wire \top.cb_syn.char_path_n[97] ;
 wire \top.cb_syn.char_path_n[98] ;
 wire \top.cb_syn.char_path_n[99] ;
 wire \top.cb_syn.char_path_n[9] ;
 wire \top.cb_syn.check_right ;
 wire \top.cb_syn.count[0] ;
 wire \top.cb_syn.count[1] ;
 wire \top.cb_syn.count[2] ;
 wire \top.cb_syn.count[3] ;
 wire \top.cb_syn.count[4] ;
 wire \top.cb_syn.count[5] ;
 wire \top.cb_syn.count[6] ;
 wire \top.cb_syn.count[7] ;
 wire \top.cb_syn.curr_index[1] ;
 wire \top.cb_syn.curr_index[2] ;
 wire \top.cb_syn.curr_index[3] ;
 wire \top.cb_syn.curr_index[4] ;
 wire \top.cb_syn.curr_index[5] ;
 wire \top.cb_syn.curr_index[6] ;
 wire \top.cb_syn.curr_index[7] ;
 wire \top.cb_syn.curr_path[127] ;
 wire \top.cb_syn.curr_state[0] ;
 wire \top.cb_syn.curr_state[1] ;
 wire \top.cb_syn.curr_state[2] ;
 wire \top.cb_syn.curr_state[4] ;
 wire \top.cb_syn.curr_state[5] ;
 wire \top.cb_syn.curr_state[8] ;
 wire \top.cb_syn.end_check ;
 wire \top.cb_syn.end_cnt[0] ;
 wire \top.cb_syn.end_cnt[1] ;
 wire \top.cb_syn.end_cnt[2] ;
 wire \top.cb_syn.end_cnt[3] ;
 wire \top.cb_syn.end_cnt[4] ;
 wire \top.cb_syn.end_cnt[5] ;
 wire \top.cb_syn.end_cnt[6] ;
 wire \top.cb_syn.end_cond ;
 wire \top.cb_syn.finished ;
 wire \top.cb_syn.h_element[46] ;
 wire \top.cb_syn.h_element[47] ;
 wire \top.cb_syn.h_element[48] ;
 wire \top.cb_syn.h_element[49] ;
 wire \top.cb_syn.h_element[50] ;
 wire \top.cb_syn.h_element[51] ;
 wire \top.cb_syn.h_element[52] ;
 wire \top.cb_syn.h_element[53] ;
 wire \top.cb_syn.h_element[54] ;
 wire \top.cb_syn.h_element[55] ;
 wire \top.cb_syn.h_element[56] ;
 wire \top.cb_syn.h_element[57] ;
 wire \top.cb_syn.h_element[58] ;
 wire \top.cb_syn.h_element[59] ;
 wire \top.cb_syn.h_element[60] ;
 wire \top.cb_syn.h_element[61] ;
 wire \top.cb_syn.h_element[62] ;
 wire \top.cb_syn.h_element[63] ;
 wire \top.cb_syn.i[0] ;
 wire \top.cb_syn.i[1] ;
 wire \top.cb_syn.i[2] ;
 wire \top.cb_syn.i[3] ;
 wire \top.cb_syn.i[4] ;
 wire \top.cb_syn.i[5] ;
 wire \top.cb_syn.i[6] ;
 wire \top.cb_syn.left ;
 wire \top.cb_syn.left_check ;
 wire \top.cb_syn.max_index[1] ;
 wire \top.cb_syn.max_index[2] ;
 wire \top.cb_syn.max_index[3] ;
 wire \top.cb_syn.max_index[4] ;
 wire \top.cb_syn.max_index[5] ;
 wire \top.cb_syn.max_index[6] ;
 wire \top.cb_syn.max_index[7] ;
 wire \top.cb_syn.num_lefts[0] ;
 wire \top.cb_syn.num_lefts[1] ;
 wire \top.cb_syn.num_lefts[2] ;
 wire \top.cb_syn.num_lefts[3] ;
 wire \top.cb_syn.num_lefts[4] ;
 wire \top.cb_syn.num_lefts[5] ;
 wire \top.cb_syn.num_lefts[6] ;
 wire \top.cb_syn.num_lefts[7] ;
 wire \top.cb_syn.pulse_first ;
 wire \top.cb_syn.pulse_first_n ;
 wire \top.cb_syn.setup ;
 wire \top.cb_syn.state8 ;
 wire \top.cb_syn.wait_cycle ;
 wire \top.cb_syn.zero_count[0] ;
 wire \top.cb_syn.zero_count[1] ;
 wire \top.cb_syn.zero_count[2] ;
 wire \top.cb_syn.zero_count[3] ;
 wire \top.cb_syn.zero_count[4] ;
 wire \top.cb_syn.zero_count[5] ;
 wire \top.cb_syn.zero_count[6] ;
 wire \top.cb_syn.zero_count[7] ;
 wire \top.cb_syn.zeroes[0] ;
 wire \top.cb_syn.zeroes[1] ;
 wire \top.cb_syn.zeroes[2] ;
 wire \top.cb_syn.zeroes[3] ;
 wire \top.cb_syn.zeroes[4] ;
 wire \top.cb_syn.zeroes[5] ;
 wire \top.cb_syn.zeroes[6] ;
 wire \top.cb_syn.zeroes[7] ;
 wire \top.compVal[0] ;
 wire \top.compVal[10] ;
 wire \top.compVal[11] ;
 wire \top.compVal[12] ;
 wire \top.compVal[13] ;
 wire \top.compVal[14] ;
 wire \top.compVal[15] ;
 wire \top.compVal[16] ;
 wire \top.compVal[17] ;
 wire \top.compVal[18] ;
 wire \top.compVal[19] ;
 wire \top.compVal[1] ;
 wire \top.compVal[20] ;
 wire \top.compVal[21] ;
 wire \top.compVal[22] ;
 wire \top.compVal[23] ;
 wire \top.compVal[24] ;
 wire \top.compVal[25] ;
 wire \top.compVal[26] ;
 wire \top.compVal[27] ;
 wire \top.compVal[28] ;
 wire \top.compVal[29] ;
 wire \top.compVal[2] ;
 wire \top.compVal[30] ;
 wire \top.compVal[31] ;
 wire \top.compVal[32] ;
 wire \top.compVal[33] ;
 wire \top.compVal[34] ;
 wire \top.compVal[35] ;
 wire \top.compVal[36] ;
 wire \top.compVal[37] ;
 wire \top.compVal[38] ;
 wire \top.compVal[39] ;
 wire \top.compVal[3] ;
 wire \top.compVal[40] ;
 wire \top.compVal[41] ;
 wire \top.compVal[42] ;
 wire \top.compVal[43] ;
 wire \top.compVal[44] ;
 wire \top.compVal[45] ;
 wire \top.compVal[4] ;
 wire \top.compVal[5] ;
 wire \top.compVal[6] ;
 wire \top.compVal[7] ;
 wire \top.compVal[8] ;
 wire \top.compVal[9] ;
 wire \top.controller.fin_FINISHED ;
 wire \top.controller.fin_FLV ;
 wire \top.controller.fin_HG ;
 wire \top.controller.fin_TRN ;
 wire \top.controller.fin_reg[1] ;
 wire \top.controller.fin_reg[2] ;
 wire \top.controller.fin_reg[3] ;
 wire \top.controller.fin_reg[4] ;
 wire \top.controller.fin_reg[5] ;
 wire \top.controller.fin_reg[6] ;
 wire \top.controller.fin_reg[7] ;
 wire \top.controller.state_reg[1] ;
 wire \top.controller.state_reg[2] ;
 wire \top.controller.state_reg[4] ;
 wire \top.controller.state_reg[5] ;
 wire \top.cw1[0] ;
 wire \top.cw1[1] ;
 wire \top.cw1[2] ;
 wire \top.cw1[3] ;
 wire \top.cw1[4] ;
 wire \top.cw1[5] ;
 wire \top.cw1[6] ;
 wire \top.cw1[7] ;
 wire \top.cw2[0] ;
 wire \top.cw2[1] ;
 wire \top.cw2[2] ;
 wire \top.cw2[3] ;
 wire \top.cw2[4] ;
 wire \top.cw2[5] ;
 wire \top.cw2[6] ;
 wire \top.cw2[7] ;
 wire \top.dut.bit_buf[0] ;
 wire \top.dut.bit_buf[10] ;
 wire \top.dut.bit_buf[11] ;
 wire \top.dut.bit_buf[12] ;
 wire \top.dut.bit_buf[13] ;
 wire \top.dut.bit_buf[1] ;
 wire \top.dut.bit_buf[2] ;
 wire \top.dut.bit_buf[3] ;
 wire \top.dut.bit_buf[4] ;
 wire \top.dut.bit_buf[5] ;
 wire \top.dut.bit_buf[6] ;
 wire \top.dut.bit_buf[7] ;
 wire \top.dut.bit_buf[8] ;
 wire \top.dut.bit_buf[9] ;
 wire \top.dut.bit_buf_next[0] ;
 wire \top.dut.bit_buf_next[10] ;
 wire \top.dut.bit_buf_next[11] ;
 wire \top.dut.bit_buf_next[12] ;
 wire \top.dut.bit_buf_next[13] ;
 wire \top.dut.bit_buf_next[1] ;
 wire \top.dut.bit_buf_next[2] ;
 wire \top.dut.bit_buf_next[3] ;
 wire \top.dut.bit_buf_next[4] ;
 wire \top.dut.bit_buf_next[5] ;
 wire \top.dut.bit_buf_next[6] ;
 wire \top.dut.bit_buf_next[7] ;
 wire \top.dut.bit_buf_next[8] ;
 wire \top.dut.bit_buf_next[9] ;
 wire \top.dut.bits_in_buf[0] ;
 wire \top.dut.bits_in_buf[1] ;
 wire \top.dut.bits_in_buf[2] ;
 wire \top.dut.bits_in_buf[3] ;
 wire \top.dut.bits_in_buf_next[0] ;
 wire \top.dut.bits_in_buf_next[1] ;
 wire \top.dut.bits_in_buf_next[2] ;
 wire \top.dut.out[0] ;
 wire \top.dut.out[1] ;
 wire \top.dut.out[2] ;
 wire \top.dut.out[3] ;
 wire \top.dut.out[4] ;
 wire \top.dut.out[5] ;
 wire \top.dut.out[6] ;
 wire \top.dut.out[7] ;
 wire \top.dut.out_valid ;
 wire \top.dut.out_valid_next ;
 wire \top.findLeastValue.alternator_timer[0] ;
 wire \top.findLeastValue.alternator_timer[1] ;
 wire \top.findLeastValue.alternator_timer[2] ;
 wire \top.findLeastValue.alternator_timer[3] ;
 wire \top.findLeastValue.histo_index[0] ;
 wire \top.findLeastValue.histo_index[1] ;
 wire \top.findLeastValue.histo_index[2] ;
 wire \top.findLeastValue.histo_index[3] ;
 wire \top.findLeastValue.histo_index[4] ;
 wire \top.findLeastValue.histo_index[5] ;
 wire \top.findLeastValue.histo_index[6] ;
 wire \top.findLeastValue.histo_index[7] ;
 wire \top.findLeastValue.histo_index[8] ;
 wire \top.findLeastValue.least1[0] ;
 wire \top.findLeastValue.least1[1] ;
 wire \top.findLeastValue.least1[2] ;
 wire \top.findLeastValue.least1[3] ;
 wire \top.findLeastValue.least1[4] ;
 wire \top.findLeastValue.least1[5] ;
 wire \top.findLeastValue.least1[6] ;
 wire \top.findLeastValue.least1[7] ;
 wire \top.findLeastValue.least1[8] ;
 wire \top.findLeastValue.least2[0] ;
 wire \top.findLeastValue.least2[1] ;
 wire \top.findLeastValue.least2[2] ;
 wire \top.findLeastValue.least2[3] ;
 wire \top.findLeastValue.least2[4] ;
 wire \top.findLeastValue.least2[5] ;
 wire \top.findLeastValue.least2[6] ;
 wire \top.findLeastValue.least2[7] ;
 wire \top.findLeastValue.least2[8] ;
 wire \top.findLeastValue.startup ;
 wire \top.findLeastValue.sum[0] ;
 wire \top.findLeastValue.sum[10] ;
 wire \top.findLeastValue.sum[11] ;
 wire \top.findLeastValue.sum[12] ;
 wire \top.findLeastValue.sum[13] ;
 wire \top.findLeastValue.sum[14] ;
 wire \top.findLeastValue.sum[15] ;
 wire \top.findLeastValue.sum[16] ;
 wire \top.findLeastValue.sum[17] ;
 wire \top.findLeastValue.sum[18] ;
 wire \top.findLeastValue.sum[19] ;
 wire \top.findLeastValue.sum[1] ;
 wire \top.findLeastValue.sum[20] ;
 wire \top.findLeastValue.sum[21] ;
 wire \top.findLeastValue.sum[22] ;
 wire \top.findLeastValue.sum[23] ;
 wire \top.findLeastValue.sum[24] ;
 wire \top.findLeastValue.sum[25] ;
 wire \top.findLeastValue.sum[26] ;
 wire \top.findLeastValue.sum[27] ;
 wire \top.findLeastValue.sum[28] ;
 wire \top.findLeastValue.sum[29] ;
 wire \top.findLeastValue.sum[2] ;
 wire \top.findLeastValue.sum[30] ;
 wire \top.findLeastValue.sum[31] ;
 wire \top.findLeastValue.sum[32] ;
 wire \top.findLeastValue.sum[33] ;
 wire \top.findLeastValue.sum[34] ;
 wire \top.findLeastValue.sum[35] ;
 wire \top.findLeastValue.sum[36] ;
 wire \top.findLeastValue.sum[37] ;
 wire \top.findLeastValue.sum[38] ;
 wire \top.findLeastValue.sum[39] ;
 wire \top.findLeastValue.sum[3] ;
 wire \top.findLeastValue.sum[40] ;
 wire \top.findLeastValue.sum[41] ;
 wire \top.findLeastValue.sum[42] ;
 wire \top.findLeastValue.sum[43] ;
 wire \top.findLeastValue.sum[44] ;
 wire \top.findLeastValue.sum[45] ;
 wire \top.findLeastValue.sum[4] ;
 wire \top.findLeastValue.sum[5] ;
 wire \top.findLeastValue.sum[6] ;
 wire \top.findLeastValue.sum[7] ;
 wire \top.findLeastValue.sum[8] ;
 wire \top.findLeastValue.sum[9] ;
 wire \top.findLeastValue.val1[0] ;
 wire \top.findLeastValue.val1[10] ;
 wire \top.findLeastValue.val1[11] ;
 wire \top.findLeastValue.val1[12] ;
 wire \top.findLeastValue.val1[13] ;
 wire \top.findLeastValue.val1[14] ;
 wire \top.findLeastValue.val1[15] ;
 wire \top.findLeastValue.val1[16] ;
 wire \top.findLeastValue.val1[17] ;
 wire \top.findLeastValue.val1[18] ;
 wire \top.findLeastValue.val1[19] ;
 wire \top.findLeastValue.val1[1] ;
 wire \top.findLeastValue.val1[20] ;
 wire \top.findLeastValue.val1[21] ;
 wire \top.findLeastValue.val1[22] ;
 wire \top.findLeastValue.val1[23] ;
 wire \top.findLeastValue.val1[24] ;
 wire \top.findLeastValue.val1[25] ;
 wire \top.findLeastValue.val1[26] ;
 wire \top.findLeastValue.val1[27] ;
 wire \top.findLeastValue.val1[28] ;
 wire \top.findLeastValue.val1[29] ;
 wire \top.findLeastValue.val1[2] ;
 wire \top.findLeastValue.val1[30] ;
 wire \top.findLeastValue.val1[31] ;
 wire \top.findLeastValue.val1[32] ;
 wire \top.findLeastValue.val1[33] ;
 wire \top.findLeastValue.val1[34] ;
 wire \top.findLeastValue.val1[35] ;
 wire \top.findLeastValue.val1[36] ;
 wire \top.findLeastValue.val1[37] ;
 wire \top.findLeastValue.val1[38] ;
 wire \top.findLeastValue.val1[39] ;
 wire \top.findLeastValue.val1[3] ;
 wire \top.findLeastValue.val1[40] ;
 wire \top.findLeastValue.val1[41] ;
 wire \top.findLeastValue.val1[42] ;
 wire \top.findLeastValue.val1[43] ;
 wire \top.findLeastValue.val1[44] ;
 wire \top.findLeastValue.val1[45] ;
 wire \top.findLeastValue.val1[46] ;
 wire \top.findLeastValue.val1[4] ;
 wire \top.findLeastValue.val1[5] ;
 wire \top.findLeastValue.val1[6] ;
 wire \top.findLeastValue.val1[7] ;
 wire \top.findLeastValue.val1[8] ;
 wire \top.findLeastValue.val1[9] ;
 wire \top.findLeastValue.val2[0] ;
 wire \top.findLeastValue.val2[10] ;
 wire \top.findLeastValue.val2[11] ;
 wire \top.findLeastValue.val2[12] ;
 wire \top.findLeastValue.val2[13] ;
 wire \top.findLeastValue.val2[14] ;
 wire \top.findLeastValue.val2[15] ;
 wire \top.findLeastValue.val2[16] ;
 wire \top.findLeastValue.val2[17] ;
 wire \top.findLeastValue.val2[18] ;
 wire \top.findLeastValue.val2[19] ;
 wire \top.findLeastValue.val2[1] ;
 wire \top.findLeastValue.val2[20] ;
 wire \top.findLeastValue.val2[21] ;
 wire \top.findLeastValue.val2[22] ;
 wire \top.findLeastValue.val2[23] ;
 wire \top.findLeastValue.val2[24] ;
 wire \top.findLeastValue.val2[25] ;
 wire \top.findLeastValue.val2[26] ;
 wire \top.findLeastValue.val2[27] ;
 wire \top.findLeastValue.val2[28] ;
 wire \top.findLeastValue.val2[29] ;
 wire \top.findLeastValue.val2[2] ;
 wire \top.findLeastValue.val2[30] ;
 wire \top.findLeastValue.val2[31] ;
 wire \top.findLeastValue.val2[32] ;
 wire \top.findLeastValue.val2[33] ;
 wire \top.findLeastValue.val2[34] ;
 wire \top.findLeastValue.val2[35] ;
 wire \top.findLeastValue.val2[36] ;
 wire \top.findLeastValue.val2[37] ;
 wire \top.findLeastValue.val2[38] ;
 wire \top.findLeastValue.val2[39] ;
 wire \top.findLeastValue.val2[3] ;
 wire \top.findLeastValue.val2[40] ;
 wire \top.findLeastValue.val2[41] ;
 wire \top.findLeastValue.val2[42] ;
 wire \top.findLeastValue.val2[43] ;
 wire \top.findLeastValue.val2[44] ;
 wire \top.findLeastValue.val2[45] ;
 wire \top.findLeastValue.val2[46] ;
 wire \top.findLeastValue.val2[4] ;
 wire \top.findLeastValue.val2[5] ;
 wire \top.findLeastValue.val2[6] ;
 wire \top.findLeastValue.val2[7] ;
 wire \top.findLeastValue.val2[8] ;
 wire \top.findLeastValue.val2[9] ;
 wire \top.findLeastValue.wipe_the_char_1 ;
 wire \top.findLeastValue.wipe_the_char_2 ;
 wire \top.hTree.closing ;
 wire \top.hTree.finish_check ;
 wire \top.hTree.node_reg[0] ;
 wire \top.hTree.node_reg[10] ;
 wire \top.hTree.node_reg[11] ;
 wire \top.hTree.node_reg[12] ;
 wire \top.hTree.node_reg[13] ;
 wire \top.hTree.node_reg[14] ;
 wire \top.hTree.node_reg[15] ;
 wire \top.hTree.node_reg[16] ;
 wire \top.hTree.node_reg[17] ;
 wire \top.hTree.node_reg[18] ;
 wire \top.hTree.node_reg[19] ;
 wire \top.hTree.node_reg[1] ;
 wire \top.hTree.node_reg[20] ;
 wire \top.hTree.node_reg[21] ;
 wire \top.hTree.node_reg[22] ;
 wire \top.hTree.node_reg[23] ;
 wire \top.hTree.node_reg[24] ;
 wire \top.hTree.node_reg[25] ;
 wire \top.hTree.node_reg[26] ;
 wire \top.hTree.node_reg[27] ;
 wire \top.hTree.node_reg[28] ;
 wire \top.hTree.node_reg[29] ;
 wire \top.hTree.node_reg[2] ;
 wire \top.hTree.node_reg[30] ;
 wire \top.hTree.node_reg[31] ;
 wire \top.hTree.node_reg[32] ;
 wire \top.hTree.node_reg[33] ;
 wire \top.hTree.node_reg[34] ;
 wire \top.hTree.node_reg[35] ;
 wire \top.hTree.node_reg[36] ;
 wire \top.hTree.node_reg[37] ;
 wire \top.hTree.node_reg[38] ;
 wire \top.hTree.node_reg[39] ;
 wire \top.hTree.node_reg[3] ;
 wire \top.hTree.node_reg[40] ;
 wire \top.hTree.node_reg[41] ;
 wire \top.hTree.node_reg[42] ;
 wire \top.hTree.node_reg[43] ;
 wire \top.hTree.node_reg[44] ;
 wire \top.hTree.node_reg[45] ;
 wire \top.hTree.node_reg[46] ;
 wire \top.hTree.node_reg[47] ;
 wire \top.hTree.node_reg[48] ;
 wire \top.hTree.node_reg[49] ;
 wire \top.hTree.node_reg[4] ;
 wire \top.hTree.node_reg[50] ;
 wire \top.hTree.node_reg[51] ;
 wire \top.hTree.node_reg[52] ;
 wire \top.hTree.node_reg[53] ;
 wire \top.hTree.node_reg[54] ;
 wire \top.hTree.node_reg[55] ;
 wire \top.hTree.node_reg[56] ;
 wire \top.hTree.node_reg[57] ;
 wire \top.hTree.node_reg[58] ;
 wire \top.hTree.node_reg[59] ;
 wire \top.hTree.node_reg[5] ;
 wire \top.hTree.node_reg[60] ;
 wire \top.hTree.node_reg[61] ;
 wire \top.hTree.node_reg[62] ;
 wire \top.hTree.node_reg[63] ;
 wire \top.hTree.node_reg[6] ;
 wire \top.hTree.node_reg[7] ;
 wire \top.hTree.node_reg[8] ;
 wire \top.hTree.node_reg[9] ;
 wire \top.hTree.nullSumIndex[0] ;
 wire \top.hTree.nullSumIndex[1] ;
 wire \top.hTree.nullSumIndex[2] ;
 wire \top.hTree.nullSumIndex[3] ;
 wire \top.hTree.nullSumIndex[4] ;
 wire \top.hTree.nullSumIndex[5] ;
 wire \top.hTree.nullSumIndex[6] ;
 wire \top.hTree.nulls[46] ;
 wire \top.hTree.nulls[47] ;
 wire \top.hTree.nulls[48] ;
 wire \top.hTree.nulls[49] ;
 wire \top.hTree.nulls[50] ;
 wire \top.hTree.nulls[51] ;
 wire \top.hTree.nulls[52] ;
 wire \top.hTree.nulls[53] ;
 wire \top.hTree.nulls[54] ;
 wire \top.hTree.nulls[55] ;
 wire \top.hTree.nulls[56] ;
 wire \top.hTree.nulls[57] ;
 wire \top.hTree.nulls[58] ;
 wire \top.hTree.nulls[59] ;
 wire \top.hTree.nulls[60] ;
 wire \top.hTree.nulls[61] ;
 wire \top.hTree.nulls[62] ;
 wire \top.hTree.nulls[63] ;
 wire \top.hTree.state[0] ;
 wire \top.hTree.state[10] ;
 wire \top.hTree.state[1] ;
 wire \top.hTree.state[2] ;
 wire \top.hTree.state[3] ;
 wire \top.hTree.state[4] ;
 wire \top.hTree.state[5] ;
 wire \top.hTree.state[6] ;
 wire \top.hTree.state[7] ;
 wire \top.hTree.state[8] ;
 wire \top.hTree.state[9] ;
 wire \top.hTree.tree_reg[0] ;
 wire \top.hTree.tree_reg[10] ;
 wire \top.hTree.tree_reg[11] ;
 wire \top.hTree.tree_reg[12] ;
 wire \top.hTree.tree_reg[13] ;
 wire \top.hTree.tree_reg[14] ;
 wire \top.hTree.tree_reg[15] ;
 wire \top.hTree.tree_reg[16] ;
 wire \top.hTree.tree_reg[17] ;
 wire \top.hTree.tree_reg[18] ;
 wire \top.hTree.tree_reg[19] ;
 wire \top.hTree.tree_reg[1] ;
 wire \top.hTree.tree_reg[20] ;
 wire \top.hTree.tree_reg[21] ;
 wire \top.hTree.tree_reg[22] ;
 wire \top.hTree.tree_reg[23] ;
 wire \top.hTree.tree_reg[24] ;
 wire \top.hTree.tree_reg[25] ;
 wire \top.hTree.tree_reg[26] ;
 wire \top.hTree.tree_reg[27] ;
 wire \top.hTree.tree_reg[28] ;
 wire \top.hTree.tree_reg[29] ;
 wire \top.hTree.tree_reg[2] ;
 wire \top.hTree.tree_reg[30] ;
 wire \top.hTree.tree_reg[31] ;
 wire \top.hTree.tree_reg[32] ;
 wire \top.hTree.tree_reg[33] ;
 wire \top.hTree.tree_reg[34] ;
 wire \top.hTree.tree_reg[35] ;
 wire \top.hTree.tree_reg[36] ;
 wire \top.hTree.tree_reg[37] ;
 wire \top.hTree.tree_reg[38] ;
 wire \top.hTree.tree_reg[39] ;
 wire \top.hTree.tree_reg[3] ;
 wire \top.hTree.tree_reg[40] ;
 wire \top.hTree.tree_reg[41] ;
 wire \top.hTree.tree_reg[42] ;
 wire \top.hTree.tree_reg[43] ;
 wire \top.hTree.tree_reg[44] ;
 wire \top.hTree.tree_reg[45] ;
 wire \top.hTree.tree_reg[46] ;
 wire \top.hTree.tree_reg[47] ;
 wire \top.hTree.tree_reg[48] ;
 wire \top.hTree.tree_reg[49] ;
 wire \top.hTree.tree_reg[4] ;
 wire \top.hTree.tree_reg[50] ;
 wire \top.hTree.tree_reg[51] ;
 wire \top.hTree.tree_reg[52] ;
 wire \top.hTree.tree_reg[53] ;
 wire \top.hTree.tree_reg[54] ;
 wire \top.hTree.tree_reg[55] ;
 wire \top.hTree.tree_reg[56] ;
 wire \top.hTree.tree_reg[57] ;
 wire \top.hTree.tree_reg[58] ;
 wire \top.hTree.tree_reg[59] ;
 wire \top.hTree.tree_reg[5] ;
 wire \top.hTree.tree_reg[60] ;
 wire \top.hTree.tree_reg[61] ;
 wire \top.hTree.tree_reg[62] ;
 wire \top.hTree.tree_reg[63] ;
 wire \top.hTree.tree_reg[6] ;
 wire \top.hTree.tree_reg[7] ;
 wire \top.hTree.tree_reg[8] ;
 wire \top.hTree.tree_reg[9] ;
 wire \top.hTree.wait_cnt ;
 wire \top.hTree.write_HT_fin ;
 wire \top.header_synthesis.bit1 ;
 wire \top.header_synthesis.char_added ;
 wire \top.header_synthesis.count[0] ;
 wire \top.header_synthesis.count[1] ;
 wire \top.header_synthesis.count[2] ;
 wire \top.header_synthesis.count[3] ;
 wire \top.header_synthesis.count[4] ;
 wire \top.header_synthesis.count[5] ;
 wire \top.header_synthesis.count[6] ;
 wire \top.header_synthesis.count[7] ;
 wire \top.header_synthesis.enable ;
 wire \top.header_synthesis.header[0] ;
 wire \top.header_synthesis.header[1] ;
 wire \top.header_synthesis.header[2] ;
 wire \top.header_synthesis.header[3] ;
 wire \top.header_synthesis.header[4] ;
 wire \top.header_synthesis.header[5] ;
 wire \top.header_synthesis.header[6] ;
 wire \top.header_synthesis.header[7] ;
 wire \top.header_synthesis.header[8] ;
 wire \top.header_synthesis.next_char_added ;
 wire \top.header_synthesis.next_enable ;
 wire \top.header_synthesis.next_header[0] ;
 wire \top.header_synthesis.next_header[1] ;
 wire \top.header_synthesis.next_header[2] ;
 wire \top.header_synthesis.next_header[3] ;
 wire \top.header_synthesis.next_header[4] ;
 wire \top.header_synthesis.next_header[5] ;
 wire \top.header_synthesis.next_header[6] ;
 wire \top.header_synthesis.next_header[7] ;
 wire \top.header_synthesis.next_header[8] ;
 wire \top.header_synthesis.next_start ;
 wire \top.header_synthesis.next_write_char_path ;
 wire \top.header_synthesis.next_write_num_lefts ;
 wire \top.header_synthesis.next_write_zeroes ;
 wire \top.header_synthesis.next_zero_count[0] ;
 wire \top.header_synthesis.next_zero_count[1] ;
 wire \top.header_synthesis.next_zero_count[2] ;
 wire \top.header_synthesis.next_zero_count[3] ;
 wire \top.header_synthesis.next_zero_count[4] ;
 wire \top.header_synthesis.next_zero_count[5] ;
 wire \top.header_synthesis.next_zero_count[6] ;
 wire \top.header_synthesis.next_zero_count[7] ;
 wire \top.header_synthesis.start ;
 wire \top.header_synthesis.write_char_path ;
 wire \top.header_synthesis.write_num_lefts ;
 wire \top.header_synthesis.write_zeroes ;
 wire \top.hist_addr[0] ;
 wire \top.hist_addr[1] ;
 wire \top.hist_addr[2] ;
 wire \top.hist_addr[3] ;
 wire \top.hist_addr[4] ;
 wire \top.hist_addr[5] ;
 wire \top.hist_addr[6] ;
 wire \top.hist_data_o[0] ;
 wire \top.hist_data_o[10] ;
 wire \top.hist_data_o[11] ;
 wire \top.hist_data_o[12] ;
 wire \top.hist_data_o[13] ;
 wire \top.hist_data_o[14] ;
 wire \top.hist_data_o[15] ;
 wire \top.hist_data_o[16] ;
 wire \top.hist_data_o[17] ;
 wire \top.hist_data_o[18] ;
 wire \top.hist_data_o[19] ;
 wire \top.hist_data_o[1] ;
 wire \top.hist_data_o[20] ;
 wire \top.hist_data_o[21] ;
 wire \top.hist_data_o[22] ;
 wire \top.hist_data_o[23] ;
 wire \top.hist_data_o[24] ;
 wire \top.hist_data_o[25] ;
 wire \top.hist_data_o[26] ;
 wire \top.hist_data_o[27] ;
 wire \top.hist_data_o[28] ;
 wire \top.hist_data_o[29] ;
 wire \top.hist_data_o[2] ;
 wire \top.hist_data_o[30] ;
 wire \top.hist_data_o[31] ;
 wire \top.hist_data_o[3] ;
 wire \top.hist_data_o[4] ;
 wire \top.hist_data_o[5] ;
 wire \top.hist_data_o[6] ;
 wire \top.hist_data_o[7] ;
 wire \top.hist_data_o[8] ;
 wire \top.hist_data_o[9] ;
 wire \top.histogram.eof_n ;
 wire \top.histogram.init ;
 wire \top.histogram.init_edge ;
 wire \top.histogram.out_of_init ;
 wire \top.histogram.sram_out[0] ;
 wire \top.histogram.sram_out[10] ;
 wire \top.histogram.sram_out[11] ;
 wire \top.histogram.sram_out[12] ;
 wire \top.histogram.sram_out[13] ;
 wire \top.histogram.sram_out[14] ;
 wire \top.histogram.sram_out[15] ;
 wire \top.histogram.sram_out[16] ;
 wire \top.histogram.sram_out[17] ;
 wire \top.histogram.sram_out[18] ;
 wire \top.histogram.sram_out[19] ;
 wire \top.histogram.sram_out[1] ;
 wire \top.histogram.sram_out[20] ;
 wire \top.histogram.sram_out[21] ;
 wire \top.histogram.sram_out[22] ;
 wire \top.histogram.sram_out[23] ;
 wire \top.histogram.sram_out[24] ;
 wire \top.histogram.sram_out[25] ;
 wire \top.histogram.sram_out[26] ;
 wire \top.histogram.sram_out[27] ;
 wire \top.histogram.sram_out[28] ;
 wire \top.histogram.sram_out[29] ;
 wire \top.histogram.sram_out[2] ;
 wire \top.histogram.sram_out[30] ;
 wire \top.histogram.sram_out[31] ;
 wire \top.histogram.sram_out[3] ;
 wire \top.histogram.sram_out[4] ;
 wire \top.histogram.sram_out[5] ;
 wire \top.histogram.sram_out[6] ;
 wire \top.histogram.sram_out[7] ;
 wire \top.histogram.sram_out[8] ;
 wire \top.histogram.sram_out[9] ;
 wire \top.histogram.state[0] ;
 wire \top.histogram.state[1] ;
 wire \top.histogram.state[2] ;
 wire \top.histogram.state[3] ;
 wire \top.histogram.state[5] ;
 wire \top.histogram.state[6] ;
 wire \top.histogram.state[7] ;
 wire \top.histogram.total[0] ;
 wire \top.histogram.total[10] ;
 wire \top.histogram.total[11] ;
 wire \top.histogram.total[12] ;
 wire \top.histogram.total[13] ;
 wire \top.histogram.total[14] ;
 wire \top.histogram.total[15] ;
 wire \top.histogram.total[16] ;
 wire \top.histogram.total[17] ;
 wire \top.histogram.total[18] ;
 wire \top.histogram.total[19] ;
 wire \top.histogram.total[1] ;
 wire \top.histogram.total[20] ;
 wire \top.histogram.total[21] ;
 wire \top.histogram.total[22] ;
 wire \top.histogram.total[23] ;
 wire \top.histogram.total[24] ;
 wire \top.histogram.total[25] ;
 wire \top.histogram.total[26] ;
 wire \top.histogram.total[27] ;
 wire \top.histogram.total[28] ;
 wire \top.histogram.total[29] ;
 wire \top.histogram.total[2] ;
 wire \top.histogram.total[30] ;
 wire \top.histogram.total[31] ;
 wire \top.histogram.total[3] ;
 wire \top.histogram.total[4] ;
 wire \top.histogram.total[5] ;
 wire \top.histogram.total[6] ;
 wire \top.histogram.total[7] ;
 wire \top.histogram.total[8] ;
 wire \top.histogram.total[9] ;
 wire \top.histogram.wr_r_en[0] ;
 wire \top.histogram.wr_r_en[1] ;
 wire \top.path[0] ;
 wire \top.path[100] ;
 wire \top.path[101] ;
 wire \top.path[102] ;
 wire \top.path[103] ;
 wire \top.path[104] ;
 wire \top.path[105] ;
 wire \top.path[106] ;
 wire \top.path[107] ;
 wire \top.path[108] ;
 wire \top.path[109] ;
 wire \top.path[10] ;
 wire \top.path[110] ;
 wire \top.path[111] ;
 wire \top.path[112] ;
 wire \top.path[113] ;
 wire \top.path[114] ;
 wire \top.path[115] ;
 wire \top.path[116] ;
 wire \top.path[117] ;
 wire \top.path[118] ;
 wire \top.path[119] ;
 wire \top.path[11] ;
 wire \top.path[120] ;
 wire \top.path[121] ;
 wire \top.path[122] ;
 wire \top.path[123] ;
 wire \top.path[124] ;
 wire \top.path[125] ;
 wire \top.path[126] ;
 wire \top.path[127] ;
 wire \top.path[12] ;
 wire \top.path[13] ;
 wire \top.path[14] ;
 wire \top.path[15] ;
 wire \top.path[16] ;
 wire \top.path[17] ;
 wire \top.path[18] ;
 wire \top.path[19] ;
 wire \top.path[1] ;
 wire \top.path[20] ;
 wire \top.path[21] ;
 wire \top.path[22] ;
 wire \top.path[23] ;
 wire \top.path[24] ;
 wire \top.path[25] ;
 wire \top.path[26] ;
 wire \top.path[27] ;
 wire \top.path[28] ;
 wire \top.path[29] ;
 wire \top.path[2] ;
 wire \top.path[30] ;
 wire \top.path[31] ;
 wire \top.path[32] ;
 wire \top.path[33] ;
 wire \top.path[34] ;
 wire \top.path[35] ;
 wire \top.path[36] ;
 wire \top.path[37] ;
 wire \top.path[38] ;
 wire \top.path[39] ;
 wire \top.path[3] ;
 wire \top.path[40] ;
 wire \top.path[41] ;
 wire \top.path[42] ;
 wire \top.path[43] ;
 wire \top.path[44] ;
 wire \top.path[45] ;
 wire \top.path[46] ;
 wire \top.path[47] ;
 wire \top.path[48] ;
 wire \top.path[49] ;
 wire \top.path[4] ;
 wire \top.path[50] ;
 wire \top.path[51] ;
 wire \top.path[52] ;
 wire \top.path[53] ;
 wire \top.path[54] ;
 wire \top.path[55] ;
 wire \top.path[56] ;
 wire \top.path[57] ;
 wire \top.path[58] ;
 wire \top.path[59] ;
 wire \top.path[5] ;
 wire \top.path[60] ;
 wire \top.path[61] ;
 wire \top.path[62] ;
 wire \top.path[63] ;
 wire \top.path[64] ;
 wire \top.path[65] ;
 wire \top.path[66] ;
 wire \top.path[67] ;
 wire \top.path[68] ;
 wire \top.path[69] ;
 wire \top.path[6] ;
 wire \top.path[70] ;
 wire \top.path[71] ;
 wire \top.path[72] ;
 wire \top.path[73] ;
 wire \top.path[74] ;
 wire \top.path[75] ;
 wire \top.path[76] ;
 wire \top.path[77] ;
 wire \top.path[78] ;
 wire \top.path[79] ;
 wire \top.path[7] ;
 wire \top.path[80] ;
 wire \top.path[81] ;
 wire \top.path[82] ;
 wire \top.path[83] ;
 wire \top.path[84] ;
 wire \top.path[85] ;
 wire \top.path[86] ;
 wire \top.path[87] ;
 wire \top.path[88] ;
 wire \top.path[89] ;
 wire \top.path[8] ;
 wire \top.path[90] ;
 wire \top.path[91] ;
 wire \top.path[92] ;
 wire \top.path[93] ;
 wire \top.path[94] ;
 wire \top.path[95] ;
 wire \top.path[96] ;
 wire \top.path[97] ;
 wire \top.path[98] ;
 wire \top.path[99] ;
 wire \top.path[9] ;
 wire \top.sram_interface.CB_read_counter ;
 wire \top.sram_interface.CB_write_counter[0] ;
 wire \top.sram_interface.CB_write_counter[1] ;
 wire \top.sram_interface.TRN_counter[0] ;
 wire \top.sram_interface.TRN_counter[1] ;
 wire \top.sram_interface.TRN_counter[2] ;
 wire \top.sram_interface.check ;
 wire \top.sram_interface.counter_HTREE[0] ;
 wire \top.sram_interface.counter_HTREE[1] ;
 wire \top.sram_interface.counter_HTREE[2] ;
 wire \top.sram_interface.counter_HTREE[3] ;
 wire \top.sram_interface.init_counter[0] ;
 wire \top.sram_interface.init_counter[10] ;
 wire \top.sram_interface.init_counter[11] ;
 wire \top.sram_interface.init_counter[12] ;
 wire \top.sram_interface.init_counter[13] ;
 wire \top.sram_interface.init_counter[14] ;
 wire \top.sram_interface.init_counter[15] ;
 wire \top.sram_interface.init_counter[16] ;
 wire \top.sram_interface.init_counter[17] ;
 wire \top.sram_interface.init_counter[18] ;
 wire \top.sram_interface.init_counter[19] ;
 wire \top.sram_interface.init_counter[1] ;
 wire \top.sram_interface.init_counter[20] ;
 wire \top.sram_interface.init_counter[21] ;
 wire \top.sram_interface.init_counter[22] ;
 wire \top.sram_interface.init_counter[23] ;
 wire \top.sram_interface.init_counter[2] ;
 wire \top.sram_interface.init_counter[3] ;
 wire \top.sram_interface.init_counter[4] ;
 wire \top.sram_interface.init_counter[5] ;
 wire \top.sram_interface.init_counter[6] ;
 wire \top.sram_interface.init_counter[7] ;
 wire \top.sram_interface.init_counter[8] ;
 wire \top.sram_interface.init_counter[9] ;
 wire \top.sram_interface.word_cnt[0] ;
 wire \top.sram_interface.word_cnt[10] ;
 wire \top.sram_interface.word_cnt[11] ;
 wire \top.sram_interface.word_cnt[12] ;
 wire \top.sram_interface.word_cnt[13] ;
 wire \top.sram_interface.word_cnt[14] ;
 wire \top.sram_interface.word_cnt[1] ;
 wire \top.sram_interface.word_cnt[2] ;
 wire \top.sram_interface.word_cnt[3] ;
 wire \top.sram_interface.word_cnt[4] ;
 wire \top.sram_interface.word_cnt[5] ;
 wire \top.sram_interface.word_cnt[6] ;
 wire \top.sram_interface.word_cnt[7] ;
 wire \top.sram_interface.word_cnt[8] ;
 wire \top.sram_interface.word_cnt[9] ;
 wire \top.sram_interface.write_HT_fin_n ;
 wire \top.sram_interface.write_counter_FLV[0] ;
 wire \top.sram_interface.write_counter_FLV[1] ;
 wire \top.sram_interface.write_counter_FLV[2] ;
 wire \top.sram_interface.zero_cnt[0] ;
 wire \top.sram_interface.zero_cnt[1] ;
 wire \top.sram_interface.zero_cnt[2] ;
 wire \top.translation.index[0] ;
 wire \top.translation.index[1] ;
 wire \top.translation.index[2] ;
 wire \top.translation.index[3] ;
 wire \top.translation.index[4] ;
 wire \top.translation.index[5] ;
 wire \top.translation.index[6] ;
 wire \top.translation.resEn ;
 wire \top.translation.totalEn ;
 wire \top.translation.writeBin ;
 wire \top.translation.writeEn ;
 wire \top.translation.write_fin ;
 wire net918;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_120_clk;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;

 sky130_fd_sc_hd__inv_2 _05287_ (.A(net441),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02404_));
 sky130_fd_sc_hd__inv_2 _05288_ (.A(net715),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02405_));
 sky130_fd_sc_hd__inv_2 _05289_ (.A(\top.compVal[45] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02406_));
 sky130_fd_sc_hd__inv_2 _05290_ (.A(\top.compVal[44] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02407_));
 sky130_fd_sc_hd__inv_2 _05291_ (.A(\top.compVal[43] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02408_));
 sky130_fd_sc_hd__inv_2 _05292_ (.A(\top.compVal[38] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02409_));
 sky130_fd_sc_hd__inv_2 _05293_ (.A(\top.compVal[37] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02410_));
 sky130_fd_sc_hd__inv_2 _05294_ (.A(\top.compVal[36] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02411_));
 sky130_fd_sc_hd__inv_2 _05295_ (.A(\top.compVal[35] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02412_));
 sky130_fd_sc_hd__inv_2 _05296_ (.A(\top.compVal[34] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02413_));
 sky130_fd_sc_hd__inv_2 _05297_ (.A(\top.compVal[33] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02414_));
 sky130_fd_sc_hd__inv_2 _05298_ (.A(\top.compVal[32] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02415_));
 sky130_fd_sc_hd__inv_2 _05299_ (.A(net481),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02416_));
 sky130_fd_sc_hd__inv_2 _05300_ (.A(net454),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02417_));
 sky130_fd_sc_hd__inv_2 _05301_ (.A(\top.hTree.write_HT_fin ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02418_));
 sky130_fd_sc_hd__inv_2 _05302_ (.A(net448),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02419_));
 sky130_fd_sc_hd__inv_2 _05303_ (.A(\top.hist_data_o[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02420_));
 sky130_fd_sc_hd__inv_2 _05304_ (.A(\top.compVal[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02421_));
 sky130_fd_sc_hd__inv_2 _05305_ (.A(\top.compVal[30] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02422_));
 sky130_fd_sc_hd__inv_2 _05306_ (.A(\top.compVal[29] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02423_));
 sky130_fd_sc_hd__inv_2 _05307_ (.A(\top.compVal[28] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02424_));
 sky130_fd_sc_hd__inv_2 _05308_ (.A(\top.compVal[27] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02425_));
 sky130_fd_sc_hd__inv_2 _05309_ (.A(\top.compVal[26] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02426_));
 sky130_fd_sc_hd__inv_2 _05310_ (.A(\top.compVal[25] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02427_));
 sky130_fd_sc_hd__inv_2 _05311_ (.A(\top.compVal[24] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02428_));
 sky130_fd_sc_hd__inv_2 _05312_ (.A(\top.compVal[23] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02429_));
 sky130_fd_sc_hd__inv_2 _05313_ (.A(\top.compVal[22] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02430_));
 sky130_fd_sc_hd__inv_2 _05314_ (.A(\top.compVal[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02431_));
 sky130_fd_sc_hd__inv_2 _05315_ (.A(\top.compVal[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02432_));
 sky130_fd_sc_hd__inv_2 _05316_ (.A(\top.compVal[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02433_));
 sky130_fd_sc_hd__inv_2 _05317_ (.A(\top.compVal[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02434_));
 sky130_fd_sc_hd__inv_2 _05318_ (.A(\top.compVal[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02435_));
 sky130_fd_sc_hd__inv_2 _05319_ (.A(\top.compVal[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02436_));
 sky130_fd_sc_hd__inv_2 _05320_ (.A(\top.compVal[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02437_));
 sky130_fd_sc_hd__inv_2 _05321_ (.A(\top.compVal[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02438_));
 sky130_fd_sc_hd__inv_2 _05322_ (.A(\top.compVal[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02439_));
 sky130_fd_sc_hd__inv_2 _05323_ (.A(\top.compVal[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02440_));
 sky130_fd_sc_hd__inv_2 _05324_ (.A(\top.compVal[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02441_));
 sky130_fd_sc_hd__inv_2 _05325_ (.A(\top.compVal[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02442_));
 sky130_fd_sc_hd__inv_2 _05326_ (.A(\top.compVal[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02443_));
 sky130_fd_sc_hd__inv_2 _05327_ (.A(\top.compVal[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02444_));
 sky130_fd_sc_hd__inv_2 _05328_ (.A(\top.compVal[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02445_));
 sky130_fd_sc_hd__inv_2 _05329_ (.A(\top.compVal[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02446_));
 sky130_fd_sc_hd__inv_2 _05330_ (.A(net981),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02447_));
 sky130_fd_sc_hd__inv_2 _05331_ (.A(\top.cb_syn.count[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02448_));
 sky130_fd_sc_hd__inv_2 _05332_ (.A(\top.cb_syn.count[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02449_));
 sky130_fd_sc_hd__inv_2 _05333_ (.A(\top.cb_syn.count[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02450_));
 sky130_fd_sc_hd__inv_2 _05334_ (.A(\top.cb_syn.count[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02451_));
 sky130_fd_sc_hd__inv_2 _05335_ (.A(\top.cb_syn.count[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02452_));
 sky130_fd_sc_hd__inv_2 _05336_ (.A(\top.cb_syn.count[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02453_));
 sky130_fd_sc_hd__inv_2 _05337_ (.A(\top.histogram.eof_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02454_));
 sky130_fd_sc_hd__inv_2 _05338_ (.A(\top.findLeastValue.val2[44] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02455_));
 sky130_fd_sc_hd__inv_2 _05339_ (.A(\top.findLeastValue.val2[42] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02456_));
 sky130_fd_sc_hd__inv_2 _05340_ (.A(\top.findLeastValue.val2[41] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02457_));
 sky130_fd_sc_hd__inv_2 _05341_ (.A(\top.findLeastValue.val2[40] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02458_));
 sky130_fd_sc_hd__inv_2 _05342_ (.A(\top.findLeastValue.val2[39] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02459_));
 sky130_fd_sc_hd__inv_2 _05343_ (.A(\top.findLeastValue.val2[37] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02460_));
 sky130_fd_sc_hd__inv_2 _05344_ (.A(\top.findLeastValue.val2[36] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02461_));
 sky130_fd_sc_hd__inv_2 _05345_ (.A(\top.findLeastValue.val2[35] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02462_));
 sky130_fd_sc_hd__inv_2 _05346_ (.A(\top.findLeastValue.val2[34] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02463_));
 sky130_fd_sc_hd__inv_2 _05347_ (.A(\top.findLeastValue.val2[33] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02464_));
 sky130_fd_sc_hd__inv_2 _05348_ (.A(\top.findLeastValue.val2[29] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02465_));
 sky130_fd_sc_hd__inv_2 _05349_ (.A(\top.findLeastValue.val2[28] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02466_));
 sky130_fd_sc_hd__inv_2 _05350_ (.A(\top.findLeastValue.val2[26] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02467_));
 sky130_fd_sc_hd__inv_2 _05351_ (.A(\top.findLeastValue.val2[24] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02468_));
 sky130_fd_sc_hd__inv_2 _05352_ (.A(\top.findLeastValue.val2[19] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02469_));
 sky130_fd_sc_hd__inv_2 _05353_ (.A(\top.findLeastValue.val2[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02470_));
 sky130_fd_sc_hd__inv_2 _05354_ (.A(\top.findLeastValue.val2[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02471_));
 sky130_fd_sc_hd__inv_2 _05355_ (.A(\top.findLeastValue.val2[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02472_));
 sky130_fd_sc_hd__inv_2 _05356_ (.A(\top.findLeastValue.val2[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02473_));
 sky130_fd_sc_hd__inv_2 _05357_ (.A(\top.findLeastValue.val2[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02474_));
 sky130_fd_sc_hd__inv_2 _05358_ (.A(\top.findLeastValue.val2[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02475_));
 sky130_fd_sc_hd__inv_2 _05359_ (.A(\top.findLeastValue.val2[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02476_));
 sky130_fd_sc_hd__inv_2 _05360_ (.A(\top.findLeastValue.val2[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02477_));
 sky130_fd_sc_hd__inv_2 _05361_ (.A(\top.findLeastValue.val2[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02478_));
 sky130_fd_sc_hd__inv_2 _05362_ (.A(\top.findLeastValue.val2[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02479_));
 sky130_fd_sc_hd__inv_2 _05363_ (.A(\top.findLeastValue.val1[44] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02480_));
 sky130_fd_sc_hd__inv_2 _05364_ (.A(\top.findLeastValue.val1[42] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02481_));
 sky130_fd_sc_hd__inv_2 _05365_ (.A(\top.findLeastValue.val1[41] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02482_));
 sky130_fd_sc_hd__inv_2 _05366_ (.A(\top.findLeastValue.val1[40] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02483_));
 sky130_fd_sc_hd__inv_2 _05367_ (.A(\top.findLeastValue.val1[39] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02484_));
 sky130_fd_sc_hd__inv_2 _05368_ (.A(\top.findLeastValue.val1[38] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02485_));
 sky130_fd_sc_hd__inv_2 _05369_ (.A(\top.findLeastValue.val1[37] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02486_));
 sky130_fd_sc_hd__inv_2 _05370_ (.A(\top.findLeastValue.val1[35] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02487_));
 sky130_fd_sc_hd__inv_2 _05371_ (.A(\top.findLeastValue.val1[33] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02488_));
 sky130_fd_sc_hd__inv_2 _05372_ (.A(\top.findLeastValue.val1[32] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02489_));
 sky130_fd_sc_hd__inv_2 _05373_ (.A(\top.findLeastValue.val1[27] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02490_));
 sky130_fd_sc_hd__inv_2 _05374_ (.A(\top.findLeastValue.val1[26] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02491_));
 sky130_fd_sc_hd__inv_2 _05375_ (.A(\top.findLeastValue.val1[21] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02492_));
 sky130_fd_sc_hd__inv_2 _05376_ (.A(\top.findLeastValue.val1[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02493_));
 sky130_fd_sc_hd__inv_2 _05377_ (.A(\top.findLeastValue.val1[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02494_));
 sky130_fd_sc_hd__inv_2 _05378_ (.A(\top.findLeastValue.val1[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02495_));
 sky130_fd_sc_hd__inv_2 _05379_ (.A(\top.findLeastValue.val1[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02496_));
 sky130_fd_sc_hd__inv_2 _05380_ (.A(\top.findLeastValue.val1[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02497_));
 sky130_fd_sc_hd__inv_2 _05381_ (.A(\top.findLeastValue.val1[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02498_));
 sky130_fd_sc_hd__inv_2 _05382_ (.A(\top.findLeastValue.wipe_the_char_2 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02499_));
 sky130_fd_sc_hd__inv_2 _05383_ (.A(\top.findLeastValue.histo_index[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02500_));
 sky130_fd_sc_hd__inv_2 _05384_ (.A(\top.findLeastValue.histo_index[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02501_));
 sky130_fd_sc_hd__inv_2 _05385_ (.A(net482),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02502_));
 sky130_fd_sc_hd__inv_2 _05386_ (.A(net483),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02503_));
 sky130_fd_sc_hd__inv_2 _05387_ (.A(\top.findLeastValue.histo_index[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02504_));
 sky130_fd_sc_hd__inv_2 _05388_ (.A(\top.cw2[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02505_));
 sky130_fd_sc_hd__inv_2 _05389_ (.A(\top.cw2[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02506_));
 sky130_fd_sc_hd__inv_2 _05390_ (.A(\top.cw2[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02507_));
 sky130_fd_sc_hd__inv_2 _05391_ (.A(\top.cw2[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02508_));
 sky130_fd_sc_hd__inv_2 _05392_ (.A(\top.cw2[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02509_));
 sky130_fd_sc_hd__inv_2 _05393_ (.A(\top.cw2[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02510_));
 sky130_fd_sc_hd__inv_2 _05394_ (.A(\top.cw2[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02511_));
 sky130_fd_sc_hd__inv_2 _05395_ (.A(\top.cw2[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02512_));
 sky130_fd_sc_hd__inv_2 _05396_ (.A(\top.cw1[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02513_));
 sky130_fd_sc_hd__inv_2 _05397_ (.A(\top.findLeastValue.least2[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02514_));
 sky130_fd_sc_hd__inv_2 _05398_ (.A(\top.findLeastValue.least2[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02515_));
 sky130_fd_sc_hd__inv_2 _05399_ (.A(\top.findLeastValue.least2[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02516_));
 sky130_fd_sc_hd__inv_2 _05400_ (.A(\top.findLeastValue.least2[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02517_));
 sky130_fd_sc_hd__inv_2 _05401_ (.A(\top.findLeastValue.least2[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02518_));
 sky130_fd_sc_hd__inv_2 _05402_ (.A(\top.findLeastValue.least2[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02519_));
 sky130_fd_sc_hd__inv_2 _05403_ (.A(\top.findLeastValue.least2[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02520_));
 sky130_fd_sc_hd__inv_2 _05404_ (.A(\top.findLeastValue.least2[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02521_));
 sky130_fd_sc_hd__inv_2 _05405_ (.A(\top.findLeastValue.least1[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02522_));
 sky130_fd_sc_hd__inv_2 _05406_ (.A(\top.findLeastValue.least1[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02523_));
 sky130_fd_sc_hd__inv_2 _05407_ (.A(\top.WorR ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02524_));
 sky130_fd_sc_hd__inv_2 _05408_ (.A(net1675),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02525_));
 sky130_fd_sc_hd__inv_2 _05409_ (.A(\top.cb_syn.zeroes[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02526_));
 sky130_fd_sc_hd__inv_2 _05410_ (.A(\top.cb_syn.zeroes[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02527_));
 sky130_fd_sc_hd__inv_2 _05411_ (.A(\top.cb_syn.zeroes[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02528_));
 sky130_fd_sc_hd__inv_2 _05412_ (.A(\top.cb_syn.zeroes[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02529_));
 sky130_fd_sc_hd__inv_2 _05413_ (.A(\top.cb_syn.zeroes[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02530_));
 sky130_fd_sc_hd__inv_2 _05414_ (.A(\top.cb_syn.zeroes[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02531_));
 sky130_fd_sc_hd__inv_2 _05415_ (.A(\top.cb_syn.zeroes[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02532_));
 sky130_fd_sc_hd__inv_2 _05416_ (.A(\top.cb_syn.zeroes[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02533_));
 sky130_fd_sc_hd__inv_2 _05417_ (.A(\top.cb_syn.cb_length[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02534_));
 sky130_fd_sc_hd__inv_2 _05418_ (.A(\top.cb_syn.cb_length[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02535_));
 sky130_fd_sc_hd__inv_2 _05419_ (.A(\top.cb_syn.char_index[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02536_));
 sky130_fd_sc_hd__inv_2 _05420_ (.A(\top.cb_syn.char_index[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02537_));
 sky130_fd_sc_hd__inv_2 _05421_ (.A(\top.cb_syn.char_path_n[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02538_));
 sky130_fd_sc_hd__inv_2 _05422_ (.A(\top.cb_syn.left_check ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02539_));
 sky130_fd_sc_hd__inv_2 _05423_ (.A(\top.cb_syn.end_cnt[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02540_));
 sky130_fd_sc_hd__inv_2 _05424_ (.A(\top.cb_syn.end_cnt[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02541_));
 sky130_fd_sc_hd__inv_2 _05425_ (.A(net496),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02542_));
 sky130_fd_sc_hd__inv_2 _05426_ (.A(net516),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02543_));
 sky130_fd_sc_hd__inv_2 _05427_ (.A(\top.header_synthesis.count[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02544_));
 sky130_fd_sc_hd__inv_2 _05428_ (.A(\top.translation.index[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02545_));
 sky130_fd_sc_hd__inv_2 _05429_ (.A(\top.translation.index[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02546_));
 sky130_fd_sc_hd__inv_2 _05430_ (.A(net503),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02547_));
 sky130_fd_sc_hd__inv_2 _05431_ (.A(net504),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02548_));
 sky130_fd_sc_hd__inv_2 _05432_ (.A(net507),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02549_));
 sky130_fd_sc_hd__inv_2 _05433_ (.A(net513),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02550_));
 sky130_fd_sc_hd__inv_2 _05434_ (.A(net550),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02551_));
 sky130_fd_sc_hd__inv_2 _05435_ (.A(\top.cb_syn.h_element[54] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02552_));
 sky130_fd_sc_hd__inv_2 _05436_ (.A(net544),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02553_));
 sky130_fd_sc_hd__inv_2 _05437_ (.A(net523),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02554_));
 sky130_fd_sc_hd__inv_2 _05438_ (.A(net463),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02555_));
 sky130_fd_sc_hd__inv_2 _05439_ (.A(\top.cb_syn.zero_count[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02556_));
 sky130_fd_sc_hd__inv_2 _05440_ (.A(\top.cb_syn.zero_count[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02557_));
 sky130_fd_sc_hd__inv_2 _05441_ (.A(\top.cb_syn.zero_count[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02558_));
 sky130_fd_sc_hd__inv_2 _05442_ (.A(\top.cb_syn.zero_count[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02559_));
 sky130_fd_sc_hd__inv_2 _05443_ (.A(net470),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02560_));
 sky130_fd_sc_hd__inv_2 _05444_ (.A(\top.dut.out_valid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02561_));
 sky130_fd_sc_hd__clkinv_4 _05445_ (.A(net455),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02562_));
 sky130_fd_sc_hd__inv_2 _05446_ (.A(net535),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02563_));
 sky130_fd_sc_hd__inv_2 _05447_ (.A(\top.sram_interface.word_cnt[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02564_));
 sky130_fd_sc_hd__inv_2 _05448_ (.A(\top.header_synthesis.enable ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02565_));
 sky130_fd_sc_hd__inv_2 _05449_ (.A(\top.header_synthesis.write_num_lefts ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02566_));
 sky130_fd_sc_hd__inv_2 _05450_ (.A(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02567_));
 sky130_fd_sc_hd__and2_1 _05451_ (.A(\top.WB.curr_state[1] ),
    .B(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02568_));
 sky130_fd_sc_hd__nand2_1 _05452_ (.A(\top.WB.curr_state[1] ),
    .B(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02569_));
 sky130_fd_sc_hd__and3_1 _05453_ (.A(net440),
    .B(\top.WB.prev_BUSY_O ),
    .C(net414),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02570_));
 sky130_fd_sc_hd__or3b_1 _05454_ (.A(net72),
    .B(net415),
    .C_N(\top.WB.prev_BUSY_O ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02571_));
 sky130_fd_sc_hd__o22a_1 _05455_ (.A1(net26),
    .A2(net414),
    .B1(net363),
    .B2(\top.WB.CPU_DAT_O[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02403_));
 sky130_fd_sc_hd__a22o_1 _05456_ (.A1(net25),
    .A2(net415),
    .B1(net364),
    .B2(\top.WB.CPU_DAT_O[30] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02402_));
 sky130_fd_sc_hd__o22a_1 _05457_ (.A1(net23),
    .A2(net413),
    .B1(net362),
    .B2(\top.WB.CPU_DAT_O[29] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02401_));
 sky130_fd_sc_hd__o22a_1 _05458_ (.A1(net22),
    .A2(net413),
    .B1(net362),
    .B2(\top.WB.CPU_DAT_O[28] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02400_));
 sky130_fd_sc_hd__o22a_1 _05459_ (.A1(net21),
    .A2(net414),
    .B1(net363),
    .B2(\top.WB.CPU_DAT_O[27] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02399_));
 sky130_fd_sc_hd__a22o_1 _05460_ (.A1(net20),
    .A2(net416),
    .B1(_02570_),
    .B2(\top.WB.CPU_DAT_O[26] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02398_));
 sky130_fd_sc_hd__o22a_1 _05461_ (.A1(net19),
    .A2(net414),
    .B1(net363),
    .B2(\top.WB.CPU_DAT_O[25] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02397_));
 sky130_fd_sc_hd__a22o_1 _05462_ (.A1(net18),
    .A2(net415),
    .B1(net364),
    .B2(\top.WB.CPU_DAT_O[24] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02396_));
 sky130_fd_sc_hd__o22a_1 _05463_ (.A1(net17),
    .A2(net414),
    .B1(net363),
    .B2(\top.WB.CPU_DAT_O[23] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02395_));
 sky130_fd_sc_hd__o22a_1 _05464_ (.A1(net16),
    .A2(net414),
    .B1(net363),
    .B2(\top.WB.CPU_DAT_O[22] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02394_));
 sky130_fd_sc_hd__a22o_1 _05465_ (.A1(net15),
    .A2(net415),
    .B1(net364),
    .B2(\top.WB.CPU_DAT_O[21] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02393_));
 sky130_fd_sc_hd__o22a_1 _05466_ (.A1(net14),
    .A2(net413),
    .B1(net362),
    .B2(\top.WB.CPU_DAT_O[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02392_));
 sky130_fd_sc_hd__a22o_1 _05467_ (.A1(net12),
    .A2(net415),
    .B1(net364),
    .B2(\top.WB.CPU_DAT_O[19] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02391_));
 sky130_fd_sc_hd__a22o_1 _05468_ (.A1(net11),
    .A2(net416),
    .B1(net364),
    .B2(\top.WB.CPU_DAT_O[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02390_));
 sky130_fd_sc_hd__a22o_1 _05469_ (.A1(net10),
    .A2(net416),
    .B1(_02570_),
    .B2(\top.WB.CPU_DAT_O[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02389_));
 sky130_fd_sc_hd__o22a_1 _05470_ (.A1(net9),
    .A2(net413),
    .B1(net363),
    .B2(\top.WB.CPU_DAT_O[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02388_));
 sky130_fd_sc_hd__o22a_1 _05471_ (.A1(net8),
    .A2(net413),
    .B1(net362),
    .B2(\top.WB.CPU_DAT_O[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02387_));
 sky130_fd_sc_hd__a22o_1 _05472_ (.A1(net7),
    .A2(net415),
    .B1(net364),
    .B2(\top.WB.CPU_DAT_O[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02386_));
 sky130_fd_sc_hd__o22a_1 _05473_ (.A1(net6),
    .A2(net413),
    .B1(net363),
    .B2(\top.WB.CPU_DAT_O[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02385_));
 sky130_fd_sc_hd__o22a_1 _05474_ (.A1(net5),
    .A2(net413),
    .B1(net362),
    .B2(\top.WB.CPU_DAT_O[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02384_));
 sky130_fd_sc_hd__o22a_1 _05475_ (.A1(net4),
    .A2(net414),
    .B1(net362),
    .B2(\top.WB.CPU_DAT_O[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02383_));
 sky130_fd_sc_hd__a22o_1 _05476_ (.A1(net3),
    .A2(net415),
    .B1(net364),
    .B2(\top.WB.CPU_DAT_O[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02382_));
 sky130_fd_sc_hd__o22a_1 _05477_ (.A1(net33),
    .A2(net413),
    .B1(net363),
    .B2(\top.WB.CPU_DAT_O[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02381_));
 sky130_fd_sc_hd__a22o_1 _05478_ (.A1(net32),
    .A2(net415),
    .B1(net364),
    .B2(\top.WB.CPU_DAT_O[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02380_));
 sky130_fd_sc_hd__o22a_1 _05479_ (.A1(net31),
    .A2(net413),
    .B1(net362),
    .B2(\top.WB.CPU_DAT_O[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02379_));
 sky130_fd_sc_hd__o22a_1 _05480_ (.A1(net30),
    .A2(net413),
    .B1(net362),
    .B2(\top.WB.CPU_DAT_O[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02378_));
 sky130_fd_sc_hd__a22o_1 _05481_ (.A1(net29),
    .A2(net415),
    .B1(net364),
    .B2(\top.WB.CPU_DAT_O[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02377_));
 sky130_fd_sc_hd__o22a_1 _05482_ (.A1(net28),
    .A2(net414),
    .B1(net362),
    .B2(\top.WB.CPU_DAT_O[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02376_));
 sky130_fd_sc_hd__a22o_1 _05483_ (.A1(net27),
    .A2(net416),
    .B1(_02570_),
    .B2(\top.WB.CPU_DAT_O[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02375_));
 sky130_fd_sc_hd__a22o_1 _05484_ (.A1(net24),
    .A2(net416),
    .B1(_02570_),
    .B2(\top.WB.CPU_DAT_O[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02374_));
 sky130_fd_sc_hd__a22o_1 _05485_ (.A1(net13),
    .A2(net415),
    .B1(net364),
    .B2(\top.WB.CPU_DAT_O[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02373_));
 sky130_fd_sc_hd__o22a_1 _05486_ (.A1(net2),
    .A2(net414),
    .B1(net362),
    .B2(\top.WB.CPU_DAT_O[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02372_));
 sky130_fd_sc_hd__nor2_1 _05487_ (.A(\top.WB.curr_state[2] ),
    .B(\top.WB.curr_state[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02572_));
 sky130_fd_sc_hd__or4_1 _05488_ (.A(net483),
    .B(net485),
    .C(net486),
    .D(\top.findLeastValue.histo_index[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02573_));
 sky130_fd_sc_hd__or2_1 _05489_ (.A(net487),
    .B(\top.findLeastValue.histo_index[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02574_));
 sky130_fd_sc_hd__or4_2 _05490_ (.A(\top.findLeastValue.histo_index[7] ),
    .B(net482),
    .C(_02573_),
    .D(_02574_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02575_));
 sky130_fd_sc_hd__nor2_2 _05491_ (.A(_02500_),
    .B(_02575_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02576_));
 sky130_fd_sc_hd__nor2_1 _05492_ (.A(_02563_),
    .B(_02576_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02577_));
 sky130_fd_sc_hd__and2_1 _05493_ (.A(net439),
    .B(net526),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02578_));
 sky130_fd_sc_hd__o2bb2a_1 _05494_ (.A1_N(\top.FLV_done ),
    .A2_N(_02576_),
    .B1(_02577_),
    .B2(net361),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02579_));
 sky130_fd_sc_hd__nor2_1 _05495_ (.A(\top.CB_read_complete ),
    .B(\top.CB_write_complete ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02580_));
 sky130_fd_sc_hd__or2_1 _05496_ (.A(\top.CB_read_complete ),
    .B(\top.CB_write_complete ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02581_));
 sky130_fd_sc_hd__or3b_2 _05497_ (.A(_02581_),
    .B(\top.cb_syn.setup ),
    .C_N(net514),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02582_));
 sky130_fd_sc_hd__a21o_1 _05498_ (.A1(net535),
    .A2(_02582_),
    .B1(\top.sram_interface.word_cnt[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02583_));
 sky130_fd_sc_hd__and2_2 _05499_ (.A(net461),
    .B(_02583_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02584_));
 sky130_fd_sc_hd__nand2_2 _05500_ (.A(net451),
    .B(net545),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02585_));
 sky130_fd_sc_hd__or2_1 _05501_ (.A(net526),
    .B(net527),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02586_));
 sky130_fd_sc_hd__nor2_1 _05502_ (.A(net537),
    .B(net527),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02587_));
 sky130_fd_sc_hd__or2_2 _05503_ (.A(net537),
    .B(net528),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02588_));
 sky130_fd_sc_hd__or2_2 _05504_ (.A(net526),
    .B(_02588_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02589_));
 sky130_fd_sc_hd__and2_1 _05505_ (.A(net451),
    .B(_02589_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02590_));
 sky130_fd_sc_hd__nand2_2 _05506_ (.A(net451),
    .B(_02589_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02591_));
 sky130_fd_sc_hd__nand2_1 _05507_ (.A(_02585_),
    .B(_02591_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02592_));
 sky130_fd_sc_hd__nor2_1 _05508_ (.A(net481),
    .B(_02417_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02593_));
 sky130_fd_sc_hd__nand2_1 _05509_ (.A(_02416_),
    .B(net453),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02594_));
 sky130_fd_sc_hd__or4b_1 _05510_ (.A(net444),
    .B(\top.histogram.wr_r_en[1] ),
    .C(_02594_),
    .D_N(\top.histogram.wr_r_en[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02595_));
 sky130_fd_sc_hd__and3_1 _05511_ (.A(net447),
    .B(\top.WorR ),
    .C(net533),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02596_));
 sky130_fd_sc_hd__a21o_1 _05512_ (.A1(net447),
    .A2(net526),
    .B1(_02596_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02597_));
 sky130_fd_sc_hd__or4b_1 _05513_ (.A(_02584_),
    .B(_02592_),
    .C(_02597_),
    .D_N(_02595_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02598_));
 sky130_fd_sc_hd__a21oi_1 _05514_ (.A1(net457),
    .A2(_02579_),
    .B1(_02598_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02599_));
 sky130_fd_sc_hd__and3_2 _05515_ (.A(net440),
    .B(\top.findLeastValue.wipe_the_char_2 ),
    .C(net527),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02600_));
 sky130_fd_sc_hd__and2_1 _05516_ (.A(\top.findLeastValue.wipe_the_char_1 ),
    .B(_02576_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02601_));
 sky130_fd_sc_hd__nand2_2 _05517_ (.A(\top.findLeastValue.wipe_the_char_1 ),
    .B(_02576_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02602_));
 sky130_fd_sc_hd__nor2_2 _05518_ (.A(_02563_),
    .B(_02602_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02603_));
 sky130_fd_sc_hd__or2_1 _05519_ (.A(_02600_),
    .B(_02603_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02604_));
 sky130_fd_sc_hd__nand2_1 _05520_ (.A(net461),
    .B(net545),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02605_));
 sky130_fd_sc_hd__nor2_1 _05521_ (.A(_02563_),
    .B(_02582_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02606_));
 sky130_fd_sc_hd__o21a_2 _05522_ (.A1(_02588_),
    .A2(net309),
    .B1(net461),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02607_));
 sky130_fd_sc_hd__a221o_1 _05523_ (.A1(net460),
    .A2(net545),
    .B1(_02604_),
    .B2(net458),
    .C1(_02607_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02608_));
 sky130_fd_sc_hd__and3_1 _05524_ (.A(net450),
    .B(_02524_),
    .C(net533),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02609_));
 sky130_fd_sc_hd__nand2_1 _05525_ (.A(net481),
    .B(net453),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02610_));
 sky130_fd_sc_hd__and2_1 _05526_ (.A(net448),
    .B(net536),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02611_));
 sky130_fd_sc_hd__a2bb2o_1 _05527_ (.A1_N(\top.sram_interface.check ),
    .A2_N(_02610_),
    .B1(\top.sram_interface.word_cnt[13] ),
    .B2(net446),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02612_));
 sky130_fd_sc_hd__or3_1 _05528_ (.A(net356),
    .B(net411),
    .C(_02612_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02613_));
 sky130_fd_sc_hd__a311o_1 _05529_ (.A1(net439),
    .A2(\top.histogram.wr_r_en[1] ),
    .A3(net360),
    .B1(_02608_),
    .C1(_02613_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02614_));
 sky130_fd_sc_hd__and2_1 _05530_ (.A(_02599_),
    .B(_02614_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02615_));
 sky130_fd_sc_hd__and3_1 _05531_ (.A(\top.WB.curr_state[0] ),
    .B(_02572_),
    .C(_02615_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02616_));
 sky130_fd_sc_hd__nor2_1 _05532_ (.A(_02599_),
    .B(_02614_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02617_));
 sky130_fd_sc_hd__or3b_1 _05533_ (.A(_02615_),
    .B(_02617_),
    .C_N(\top.WB.curr_state[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02618_));
 sky130_fd_sc_hd__or3b_2 _05534_ (.A(_02567_),
    .B(_02572_),
    .C_N(_02618_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02619_));
 sky130_fd_sc_hd__a31o_1 _05535_ (.A1(\top.WB.curr_state[0] ),
    .A2(_02572_),
    .A3(_02617_),
    .B1(net213),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02620_));
 sky130_fd_sc_hd__and2b_2 _05536_ (.A_N(net207),
    .B(_02619_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02621_));
 sky130_fd_sc_hd__a21o_1 _05537_ (.A1(net1026),
    .A2(net169),
    .B1(net211),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02371_));
 sky130_fd_sc_hd__a21o_1 _05538_ (.A1(net441),
    .A2(_02619_),
    .B1(net207),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02370_));
 sky130_fd_sc_hd__a22o_1 _05539_ (.A1(\top.cb_syn.char_path[31] ),
    .A2(net546),
    .B1(net538),
    .B2(\top.cb_syn.char_path[95] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02622_));
 sky130_fd_sc_hd__a22o_1 _05540_ (.A1(\top.cb_syn.char_path[63] ),
    .A2(net528),
    .B1(net309),
    .B2(\top.cb_syn.char_path[127] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02623_));
 sky130_fd_sc_hd__o21a_1 _05541_ (.A1(_02622_),
    .A2(_02623_),
    .B1(net465),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02624_));
 sky130_fd_sc_hd__a22o_1 _05542_ (.A1(\top.histogram.sram_out[31] ),
    .A2(net360),
    .B1(net411),
    .B2(\top.hTree.node_reg[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02625_));
 sky130_fd_sc_hd__a211o_1 _05543_ (.A1(\top.hTree.node_reg[63] ),
    .A2(net356),
    .B1(_02624_),
    .C1(_02625_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02626_));
 sky130_fd_sc_hd__a22o_1 _05544_ (.A1(net97),
    .A2(net167),
    .B1(_02626_),
    .B2(net213),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02369_));
 sky130_fd_sc_hd__a22o_1 _05545_ (.A1(\top.cb_syn.char_path[30] ),
    .A2(net546),
    .B1(net538),
    .B2(\top.cb_syn.char_path[94] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02627_));
 sky130_fd_sc_hd__a22o_1 _05546_ (.A1(\top.cb_syn.char_path[62] ),
    .A2(net528),
    .B1(net309),
    .B2(\top.cb_syn.char_path[126] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02628_));
 sky130_fd_sc_hd__o21a_1 _05547_ (.A1(_02627_),
    .A2(_02628_),
    .B1(net465),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02629_));
 sky130_fd_sc_hd__a22o_1 _05548_ (.A1(\top.histogram.sram_out[30] ),
    .A2(net360),
    .B1(net411),
    .B2(\top.hTree.node_reg[30] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02630_));
 sky130_fd_sc_hd__a211o_1 _05549_ (.A1(\top.hTree.node_reg[62] ),
    .A2(net356),
    .B1(_02629_),
    .C1(_02630_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02631_));
 sky130_fd_sc_hd__a22o_1 _05550_ (.A1(net1796),
    .A2(net166),
    .B1(_02631_),
    .B2(net213),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02368_));
 sky130_fd_sc_hd__a22o_1 _05551_ (.A1(\top.cb_syn.char_path[93] ),
    .A2(net537),
    .B1(net528),
    .B2(\top.cb_syn.char_path[61] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02632_));
 sky130_fd_sc_hd__a22o_1 _05552_ (.A1(\top.cb_syn.char_path[29] ),
    .A2(net546),
    .B1(net309),
    .B2(\top.cb_syn.char_path[125] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02633_));
 sky130_fd_sc_hd__o21a_1 _05553_ (.A1(_02632_),
    .A2(_02633_),
    .B1(net465),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02634_));
 sky130_fd_sc_hd__a22o_1 _05554_ (.A1(\top.histogram.sram_out[29] ),
    .A2(net360),
    .B1(net411),
    .B2(\top.hTree.node_reg[29] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02635_));
 sky130_fd_sc_hd__a211o_1 _05555_ (.A1(\top.hTree.node_reg[61] ),
    .A2(net356),
    .B1(_02634_),
    .C1(_02635_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02636_));
 sky130_fd_sc_hd__a22o_1 _05556_ (.A1(net1777),
    .A2(net167),
    .B1(_02636_),
    .B2(net213),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02367_));
 sky130_fd_sc_hd__a22o_1 _05557_ (.A1(\top.cb_syn.char_path[28] ),
    .A2(net546),
    .B1(net537),
    .B2(\top.cb_syn.char_path[92] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02637_));
 sky130_fd_sc_hd__a22o_1 _05558_ (.A1(\top.cb_syn.char_path[60] ),
    .A2(net528),
    .B1(net309),
    .B2(\top.cb_syn.char_path[124] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02638_));
 sky130_fd_sc_hd__o21a_1 _05559_ (.A1(_02637_),
    .A2(_02638_),
    .B1(net465),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02639_));
 sky130_fd_sc_hd__a22o_1 _05560_ (.A1(\top.histogram.sram_out[28] ),
    .A2(net360),
    .B1(net411),
    .B2(\top.hTree.node_reg[28] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02640_));
 sky130_fd_sc_hd__a211o_1 _05561_ (.A1(net1799),
    .A2(net354),
    .B1(_02639_),
    .C1(_02640_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02641_));
 sky130_fd_sc_hd__a22o_1 _05562_ (.A1(net93),
    .A2(net171),
    .B1(_02641_),
    .B2(net213),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02366_));
 sky130_fd_sc_hd__a22o_1 _05563_ (.A1(\top.cb_syn.char_path[91] ),
    .A2(net537),
    .B1(net532),
    .B2(\top.cb_syn.char_path[59] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02642_));
 sky130_fd_sc_hd__a22o_1 _05564_ (.A1(\top.cb_syn.char_path[27] ),
    .A2(\top.sram_interface.word_cnt[0] ),
    .B1(net309),
    .B2(\top.cb_syn.char_path[123] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02643_));
 sky130_fd_sc_hd__o21a_1 _05565_ (.A1(_02642_),
    .A2(_02643_),
    .B1(net465),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02644_));
 sky130_fd_sc_hd__a22o_1 _05566_ (.A1(\top.hTree.node_reg[59] ),
    .A2(net354),
    .B1(net410),
    .B2(\top.hTree.node_reg[27] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02645_));
 sky130_fd_sc_hd__a211o_1 _05567_ (.A1(\top.histogram.sram_out[27] ),
    .A2(net359),
    .B1(_02644_),
    .C1(_02645_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02646_));
 sky130_fd_sc_hd__a22o_1 _05568_ (.A1(net1460),
    .A2(net170),
    .B1(_02646_),
    .B2(net209),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02365_));
 sky130_fd_sc_hd__a22o_1 _05569_ (.A1(\top.cb_syn.char_path[26] ),
    .A2(net546),
    .B1(net537),
    .B2(\top.cb_syn.char_path[90] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02647_));
 sky130_fd_sc_hd__a22o_1 _05570_ (.A1(\top.cb_syn.char_path[58] ),
    .A2(net532),
    .B1(net309),
    .B2(\top.cb_syn.char_path[122] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02648_));
 sky130_fd_sc_hd__or2_1 _05571_ (.A(_02647_),
    .B(_02648_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02649_));
 sky130_fd_sc_hd__a22o_1 _05572_ (.A1(\top.histogram.sram_out[26] ),
    .A2(net359),
    .B1(_02649_),
    .B2(net467),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02650_));
 sky130_fd_sc_hd__a221o_1 _05573_ (.A1(\top.hTree.node_reg[58] ),
    .A2(net354),
    .B1(net410),
    .B2(\top.hTree.node_reg[26] ),
    .C1(_02650_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02651_));
 sky130_fd_sc_hd__a22o_1 _05574_ (.A1(net1421),
    .A2(net168),
    .B1(_02651_),
    .B2(net210),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02364_));
 sky130_fd_sc_hd__a22o_1 _05575_ (.A1(\top.cb_syn.char_path[89] ),
    .A2(net537),
    .B1(net532),
    .B2(\top.cb_syn.char_path[57] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02652_));
 sky130_fd_sc_hd__a22o_1 _05576_ (.A1(\top.cb_syn.char_path[25] ),
    .A2(net546),
    .B1(net312),
    .B2(\top.cb_syn.char_path[121] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02653_));
 sky130_fd_sc_hd__o21a_1 _05577_ (.A1(_02652_),
    .A2(_02653_),
    .B1(net466),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02654_));
 sky130_fd_sc_hd__a22o_1 _05578_ (.A1(\top.histogram.sram_out[25] ),
    .A2(net359),
    .B1(net354),
    .B2(\top.hTree.node_reg[57] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02655_));
 sky130_fd_sc_hd__a211o_1 _05579_ (.A1(\top.hTree.node_reg[25] ),
    .A2(net410),
    .B1(_02654_),
    .C1(_02655_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02656_));
 sky130_fd_sc_hd__a22o_1 _05580_ (.A1(net1447),
    .A2(net168),
    .B1(_02656_),
    .B2(net210),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02363_));
 sky130_fd_sc_hd__a22o_1 _05581_ (.A1(\top.cb_syn.char_path[24] ),
    .A2(\top.sram_interface.word_cnt[0] ),
    .B1(net538),
    .B2(\top.cb_syn.char_path[88] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02657_));
 sky130_fd_sc_hd__a22o_1 _05582_ (.A1(\top.cb_syn.char_path[56] ),
    .A2(net528),
    .B1(net312),
    .B2(\top.cb_syn.char_path[120] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02658_));
 sky130_fd_sc_hd__o21a_1 _05583_ (.A1(_02657_),
    .A2(_02658_),
    .B1(net465),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02659_));
 sky130_fd_sc_hd__a22o_1 _05584_ (.A1(\top.histogram.sram_out[24] ),
    .A2(net359),
    .B1(net410),
    .B2(\top.hTree.node_reg[24] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02660_));
 sky130_fd_sc_hd__a211o_1 _05585_ (.A1(net1019),
    .A2(net354),
    .B1(_02659_),
    .C1(_02660_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02661_));
 sky130_fd_sc_hd__a22o_1 _05586_ (.A1(net89),
    .A2(net171),
    .B1(_02661_),
    .B2(net212),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02362_));
 sky130_fd_sc_hd__a22o_1 _05587_ (.A1(\top.cb_syn.char_path[23] ),
    .A2(net548),
    .B1(net538),
    .B2(\top.cb_syn.char_path[87] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02662_));
 sky130_fd_sc_hd__a22o_1 _05588_ (.A1(\top.cb_syn.char_path[55] ),
    .A2(net530),
    .B1(net311),
    .B2(\top.cb_syn.char_path[119] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02663_));
 sky130_fd_sc_hd__o21a_1 _05589_ (.A1(_02662_),
    .A2(_02663_),
    .B1(net467),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02664_));
 sky130_fd_sc_hd__a22o_1 _05590_ (.A1(\top.histogram.sram_out[23] ),
    .A2(net359),
    .B1(net354),
    .B2(\top.hTree.node_reg[55] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02665_));
 sky130_fd_sc_hd__a211o_1 _05591_ (.A1(\top.hTree.node_reg[23] ),
    .A2(net410),
    .B1(_02664_),
    .C1(_02665_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02666_));
 sky130_fd_sc_hd__a22o_1 _05592_ (.A1(net1211),
    .A2(net168),
    .B1(_02666_),
    .B2(net210),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02361_));
 sky130_fd_sc_hd__a22o_1 _05593_ (.A1(\top.cb_syn.char_path[22] ),
    .A2(net548),
    .B1(net539),
    .B2(\top.cb_syn.char_path[86] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02667_));
 sky130_fd_sc_hd__a22o_1 _05594_ (.A1(\top.cb_syn.char_path[54] ),
    .A2(net530),
    .B1(net311),
    .B2(\top.cb_syn.char_path[118] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02668_));
 sky130_fd_sc_hd__o21a_1 _05595_ (.A1(_02667_),
    .A2(_02668_),
    .B1(net467),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02669_));
 sky130_fd_sc_hd__a22o_1 _05596_ (.A1(\top.histogram.sram_out[22] ),
    .A2(net359),
    .B1(net354),
    .B2(\top.hTree.node_reg[54] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02670_));
 sky130_fd_sc_hd__a211o_1 _05597_ (.A1(\top.hTree.node_reg[22] ),
    .A2(net410),
    .B1(_02669_),
    .C1(_02670_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02671_));
 sky130_fd_sc_hd__a22o_1 _05598_ (.A1(net1169),
    .A2(net168),
    .B1(_02671_),
    .B2(net210),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02360_));
 sky130_fd_sc_hd__a22o_1 _05599_ (.A1(\top.cb_syn.char_path[21] ),
    .A2(net548),
    .B1(net539),
    .B2(\top.cb_syn.char_path[85] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02672_));
 sky130_fd_sc_hd__a22o_1 _05600_ (.A1(\top.cb_syn.char_path[53] ),
    .A2(net530),
    .B1(net311),
    .B2(\top.cb_syn.char_path[117] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02673_));
 sky130_fd_sc_hd__o21a_1 _05601_ (.A1(_02672_),
    .A2(_02673_),
    .B1(net467),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02674_));
 sky130_fd_sc_hd__a22o_1 _05602_ (.A1(\top.histogram.sram_out[21] ),
    .A2(net359),
    .B1(net410),
    .B2(\top.hTree.node_reg[21] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02675_));
 sky130_fd_sc_hd__a211o_1 _05603_ (.A1(\top.hTree.node_reg[53] ),
    .A2(net354),
    .B1(_02674_),
    .C1(_02675_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02676_));
 sky130_fd_sc_hd__a22o_1 _05604_ (.A1(net1484),
    .A2(net169),
    .B1(_02676_),
    .B2(net211),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02359_));
 sky130_fd_sc_hd__a22o_1 _05605_ (.A1(\top.cb_syn.char_path[20] ),
    .A2(net548),
    .B1(net539),
    .B2(\top.cb_syn.char_path[84] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02677_));
 sky130_fd_sc_hd__a22o_1 _05606_ (.A1(\top.cb_syn.char_path[52] ),
    .A2(net530),
    .B1(net311),
    .B2(\top.cb_syn.char_path[116] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02678_));
 sky130_fd_sc_hd__o21a_1 _05607_ (.A1(_02677_),
    .A2(_02678_),
    .B1(net467),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02679_));
 sky130_fd_sc_hd__a22o_1 _05608_ (.A1(\top.histogram.sram_out[20] ),
    .A2(net359),
    .B1(net410),
    .B2(\top.hTree.node_reg[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02680_));
 sky130_fd_sc_hd__a211o_1 _05609_ (.A1(\top.hTree.node_reg[52] ),
    .A2(net354),
    .B1(_02679_),
    .C1(_02680_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02681_));
 sky130_fd_sc_hd__a22o_1 _05610_ (.A1(net1477),
    .A2(net169),
    .B1(_02681_),
    .B2(net211),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02358_));
 sky130_fd_sc_hd__a22o_1 _05611_ (.A1(\top.cb_syn.char_path[19] ),
    .A2(net548),
    .B1(net539),
    .B2(\top.cb_syn.char_path[83] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02682_));
 sky130_fd_sc_hd__a22o_1 _05612_ (.A1(\top.cb_syn.char_path[51] ),
    .A2(net530),
    .B1(net311),
    .B2(\top.cb_syn.char_path[115] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02683_));
 sky130_fd_sc_hd__o21a_1 _05613_ (.A1(_02682_),
    .A2(_02683_),
    .B1(net467),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02684_));
 sky130_fd_sc_hd__a22o_1 _05614_ (.A1(\top.histogram.sram_out[19] ),
    .A2(net359),
    .B1(net410),
    .B2(\top.hTree.node_reg[19] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02685_));
 sky130_fd_sc_hd__a211o_1 _05615_ (.A1(\top.hTree.node_reg[51] ),
    .A2(net354),
    .B1(_02684_),
    .C1(_02685_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02686_));
 sky130_fd_sc_hd__a22o_1 _05616_ (.A1(net1365),
    .A2(net171),
    .B1(_02686_),
    .B2(net211),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02357_));
 sky130_fd_sc_hd__a22o_1 _05617_ (.A1(\top.cb_syn.char_path[18] ),
    .A2(net548),
    .B1(net539),
    .B2(\top.cb_syn.char_path[82] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02687_));
 sky130_fd_sc_hd__a22o_1 _05618_ (.A1(\top.cb_syn.char_path[50] ),
    .A2(net530),
    .B1(net311),
    .B2(\top.cb_syn.char_path[114] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02688_));
 sky130_fd_sc_hd__o21a_1 _05619_ (.A1(_02687_),
    .A2(_02688_),
    .B1(net467),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02689_));
 sky130_fd_sc_hd__a22o_1 _05620_ (.A1(\top.histogram.sram_out[18] ),
    .A2(net358),
    .B1(net410),
    .B2(\top.hTree.node_reg[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02690_));
 sky130_fd_sc_hd__a211o_1 _05621_ (.A1(\top.hTree.node_reg[50] ),
    .A2(net355),
    .B1(_02689_),
    .C1(_02690_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02691_));
 sky130_fd_sc_hd__a22o_1 _05622_ (.A1(net1452),
    .A2(net169),
    .B1(_02691_),
    .B2(net210),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02356_));
 sky130_fd_sc_hd__a22o_1 _05623_ (.A1(\top.cb_syn.char_path[17] ),
    .A2(net547),
    .B1(net539),
    .B2(\top.cb_syn.char_path[81] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02692_));
 sky130_fd_sc_hd__a22o_1 _05624_ (.A1(\top.cb_syn.char_path[49] ),
    .A2(net530),
    .B1(net311),
    .B2(\top.cb_syn.char_path[113] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02693_));
 sky130_fd_sc_hd__o21a_1 _05625_ (.A1(_02692_),
    .A2(_02693_),
    .B1(net468),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02694_));
 sky130_fd_sc_hd__a22o_1 _05626_ (.A1(\top.histogram.sram_out[17] ),
    .A2(net358),
    .B1(net355),
    .B2(\top.hTree.node_reg[49] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02695_));
 sky130_fd_sc_hd__a211o_1 _05627_ (.A1(\top.hTree.node_reg[17] ),
    .A2(net409),
    .B1(_02694_),
    .C1(_02695_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02696_));
 sky130_fd_sc_hd__a22o_1 _05628_ (.A1(net1196),
    .A2(net169),
    .B1(_02696_),
    .B2(net210),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02355_));
 sky130_fd_sc_hd__a22o_1 _05629_ (.A1(\top.cb_syn.char_path[16] ),
    .A2(net547),
    .B1(net540),
    .B2(\top.cb_syn.char_path[80] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02697_));
 sky130_fd_sc_hd__a22o_1 _05630_ (.A1(\top.cb_syn.char_path[48] ),
    .A2(net531),
    .B1(net310),
    .B2(\top.cb_syn.char_path[112] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02698_));
 sky130_fd_sc_hd__o21a_1 _05631_ (.A1(_02697_),
    .A2(_02698_),
    .B1(net468),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02699_));
 sky130_fd_sc_hd__a22o_1 _05632_ (.A1(\top.histogram.sram_out[16] ),
    .A2(net358),
    .B1(net355),
    .B2(\top.hTree.node_reg[48] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02700_));
 sky130_fd_sc_hd__a211o_1 _05633_ (.A1(\top.hTree.node_reg[16] ),
    .A2(net409),
    .B1(_02699_),
    .C1(_02700_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02701_));
 sky130_fd_sc_hd__a22o_1 _05634_ (.A1(net1383),
    .A2(net168),
    .B1(_02701_),
    .B2(net210),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02354_));
 sky130_fd_sc_hd__a22o_1 _05635_ (.A1(\top.cb_syn.char_path[15] ),
    .A2(net549),
    .B1(net540),
    .B2(\top.cb_syn.char_path[79] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02702_));
 sky130_fd_sc_hd__a22o_1 _05636_ (.A1(\top.cb_syn.char_path[47] ),
    .A2(net531),
    .B1(net312),
    .B2(\top.cb_syn.char_path[111] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02703_));
 sky130_fd_sc_hd__o21a_1 _05637_ (.A1(_02702_),
    .A2(_02703_),
    .B1(net468),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02704_));
 sky130_fd_sc_hd__a22o_1 _05638_ (.A1(\top.histogram.sram_out[15] ),
    .A2(net358),
    .B1(net409),
    .B2(\top.hTree.node_reg[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02705_));
 sky130_fd_sc_hd__a211o_1 _05639_ (.A1(\top.hTree.node_reg[47] ),
    .A2(net355),
    .B1(_02704_),
    .C1(_02705_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02706_));
 sky130_fd_sc_hd__a22o_1 _05640_ (.A1(net1359),
    .A2(net171),
    .B1(_02706_),
    .B2(net211),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02353_));
 sky130_fd_sc_hd__a22o_1 _05641_ (.A1(\top.cb_syn.char_path[78] ),
    .A2(net540),
    .B1(net531),
    .B2(\top.cb_syn.char_path[46] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02707_));
 sky130_fd_sc_hd__a22o_1 _05642_ (.A1(\top.cb_syn.char_path[14] ),
    .A2(net547),
    .B1(net312),
    .B2(\top.cb_syn.char_path[110] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02708_));
 sky130_fd_sc_hd__o21a_1 _05643_ (.A1(_02707_),
    .A2(_02708_),
    .B1(net468),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02709_));
 sky130_fd_sc_hd__a22o_1 _05644_ (.A1(\top.histogram.sram_out[14] ),
    .A2(net358),
    .B1(net409),
    .B2(\top.hTree.node_reg[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02710_));
 sky130_fd_sc_hd__a211o_1 _05645_ (.A1(\top.hTree.node_reg[46] ),
    .A2(net355),
    .B1(_02709_),
    .C1(_02710_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02711_));
 sky130_fd_sc_hd__a22o_1 _05646_ (.A1(net1316),
    .A2(net171),
    .B1(_02711_),
    .B2(net211),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02352_));
 sky130_fd_sc_hd__a22o_1 _05647_ (.A1(\top.cb_syn.char_path[13] ),
    .A2(net547),
    .B1(net540),
    .B2(\top.cb_syn.char_path[77] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02712_));
 sky130_fd_sc_hd__a22o_1 _05648_ (.A1(\top.cb_syn.char_path[45] ),
    .A2(net531),
    .B1(net310),
    .B2(\top.cb_syn.char_path[109] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02713_));
 sky130_fd_sc_hd__or2_1 _05649_ (.A(_02712_),
    .B(_02713_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02714_));
 sky130_fd_sc_hd__and2_1 _05650_ (.A(_02418_),
    .B(net356),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02715_));
 sky130_fd_sc_hd__a22o_1 _05651_ (.A1(net467),
    .A2(_02714_),
    .B1(net307),
    .B2(\top.hTree.node_reg[45] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02716_));
 sky130_fd_sc_hd__a221o_1 _05652_ (.A1(\top.histogram.sram_out[13] ),
    .A2(net358),
    .B1(net409),
    .B2(\top.hTree.node_reg[13] ),
    .C1(_02716_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02717_));
 sky130_fd_sc_hd__a22o_1 _05653_ (.A1(net1530),
    .A2(net168),
    .B1(_02717_),
    .B2(net210),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02351_));
 sky130_fd_sc_hd__a22o_1 _05654_ (.A1(\top.cb_syn.char_path[76] ),
    .A2(net540),
    .B1(net529),
    .B2(\top.cb_syn.char_path[44] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02718_));
 sky130_fd_sc_hd__a22o_1 _05655_ (.A1(\top.cb_syn.char_path[12] ),
    .A2(net547),
    .B1(net310),
    .B2(\top.cb_syn.char_path[108] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02719_));
 sky130_fd_sc_hd__or2_1 _05656_ (.A(_02718_),
    .B(_02719_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02720_));
 sky130_fd_sc_hd__a22o_1 _05657_ (.A1(\top.hTree.node_reg[44] ),
    .A2(net307),
    .B1(_02720_),
    .B2(net467),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02721_));
 sky130_fd_sc_hd__a221o_1 _05658_ (.A1(\top.histogram.sram_out[12] ),
    .A2(net358),
    .B1(net409),
    .B2(\top.hTree.node_reg[12] ),
    .C1(_02721_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02722_));
 sky130_fd_sc_hd__a22o_1 _05659_ (.A1(net1462),
    .A2(net168),
    .B1(_02722_),
    .B2(net210),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02350_));
 sky130_fd_sc_hd__a22o_1 _05660_ (.A1(\top.cb_syn.char_path[11] ),
    .A2(net547),
    .B1(net539),
    .B2(\top.cb_syn.char_path[75] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02723_));
 sky130_fd_sc_hd__a22o_1 _05661_ (.A1(\top.cb_syn.char_path[43] ),
    .A2(net529),
    .B1(net310),
    .B2(\top.cb_syn.char_path[107] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02724_));
 sky130_fd_sc_hd__or2_1 _05662_ (.A(_02723_),
    .B(_02724_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02725_));
 sky130_fd_sc_hd__a22o_1 _05663_ (.A1(\top.hTree.node_reg[43] ),
    .A2(net308),
    .B1(_02725_),
    .B2(net469),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02726_));
 sky130_fd_sc_hd__a221o_1 _05664_ (.A1(\top.histogram.sram_out[11] ),
    .A2(net357),
    .B1(net408),
    .B2(\top.hTree.node_reg[11] ),
    .C1(_02726_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02727_));
 sky130_fd_sc_hd__a22o_1 _05665_ (.A1(net1307),
    .A2(net168),
    .B1(_02727_),
    .B2(net210),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02349_));
 sky130_fd_sc_hd__a22o_1 _05666_ (.A1(\top.cb_syn.char_path[74] ),
    .A2(net540),
    .B1(net529),
    .B2(\top.cb_syn.char_path[42] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02728_));
 sky130_fd_sc_hd__a22o_1 _05667_ (.A1(\top.cb_syn.char_path[10] ),
    .A2(net547),
    .B1(net310),
    .B2(\top.cb_syn.char_path[106] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02729_));
 sky130_fd_sc_hd__o21a_1 _05668_ (.A1(_02728_),
    .A2(_02729_),
    .B1(net468),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02730_));
 sky130_fd_sc_hd__a22o_1 _05669_ (.A1(\top.histogram.sram_out[10] ),
    .A2(net357),
    .B1(net408),
    .B2(\top.hTree.node_reg[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02731_));
 sky130_fd_sc_hd__a211o_1 _05670_ (.A1(\top.hTree.node_reg[42] ),
    .A2(net307),
    .B1(_02730_),
    .C1(_02731_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02732_));
 sky130_fd_sc_hd__a22o_1 _05671_ (.A1(net1411),
    .A2(net168),
    .B1(_02732_),
    .B2(net209),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02348_));
 sky130_fd_sc_hd__a22o_1 _05672_ (.A1(\top.cb_syn.char_path[9] ),
    .A2(net547),
    .B1(net540),
    .B2(\top.cb_syn.char_path[73] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02733_));
 sky130_fd_sc_hd__a22o_1 _05673_ (.A1(\top.cb_syn.char_path[41] ),
    .A2(net529),
    .B1(net312),
    .B2(\top.cb_syn.char_path[105] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02734_));
 sky130_fd_sc_hd__or2_1 _05674_ (.A(_02733_),
    .B(_02734_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02735_));
 sky130_fd_sc_hd__a22o_1 _05675_ (.A1(\top.hTree.node_reg[41] ),
    .A2(net308),
    .B1(_02735_),
    .B2(net469),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02736_));
 sky130_fd_sc_hd__a221o_1 _05676_ (.A1(\top.histogram.sram_out[9] ),
    .A2(net357),
    .B1(net408),
    .B2(\top.hTree.node_reg[9] ),
    .C1(_02736_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02737_));
 sky130_fd_sc_hd__a22o_1 _05677_ (.A1(net1469),
    .A2(net168),
    .B1(_02737_),
    .B2(net209),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02347_));
 sky130_fd_sc_hd__a22o_1 _05678_ (.A1(\top.cb_syn.char_path[8] ),
    .A2(net547),
    .B1(net540),
    .B2(\top.cb_syn.char_path[72] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02738_));
 sky130_fd_sc_hd__a22o_1 _05679_ (.A1(\top.cb_syn.char_path[40] ),
    .A2(net529),
    .B1(net312),
    .B2(\top.cb_syn.char_path[104] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02739_));
 sky130_fd_sc_hd__or2_1 _05680_ (.A(_02738_),
    .B(_02739_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02740_));
 sky130_fd_sc_hd__a22o_1 _05681_ (.A1(\top.hTree.node_reg[40] ),
    .A2(net308),
    .B1(_02740_),
    .B2(net468),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02741_));
 sky130_fd_sc_hd__a221o_1 _05682_ (.A1(\top.histogram.sram_out[8] ),
    .A2(net358),
    .B1(net409),
    .B2(\top.hTree.node_reg[8] ),
    .C1(_02741_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02742_));
 sky130_fd_sc_hd__a22o_1 _05683_ (.A1(net1397),
    .A2(net169),
    .B1(_02742_),
    .B2(net211),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02346_));
 sky130_fd_sc_hd__a22o_1 _05684_ (.A1(\top.cb_syn.char_path[7] ),
    .A2(net547),
    .B1(net540),
    .B2(\top.cb_syn.char_path[71] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02743_));
 sky130_fd_sc_hd__a22o_1 _05685_ (.A1(\top.cb_syn.char_path[39] ),
    .A2(net529),
    .B1(net310),
    .B2(\top.cb_syn.char_path[103] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02744_));
 sky130_fd_sc_hd__o21a_1 _05686_ (.A1(_02743_),
    .A2(_02744_),
    .B1(net468),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02745_));
 sky130_fd_sc_hd__a22o_1 _05687_ (.A1(\top.histogram.sram_out[7] ),
    .A2(net357),
    .B1(net408),
    .B2(\top.hTree.node_reg[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02746_));
 sky130_fd_sc_hd__a211o_1 _05688_ (.A1(\top.hTree.node_reg[39] ),
    .A2(net307),
    .B1(_02745_),
    .C1(_02746_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02747_));
 sky130_fd_sc_hd__a22o_1 _05689_ (.A1(net1282),
    .A2(net170),
    .B1(_02747_),
    .B2(net209),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02345_));
 sky130_fd_sc_hd__a22o_1 _05690_ (.A1(\top.cb_syn.char_path[6] ),
    .A2(net549),
    .B1(net541),
    .B2(\top.cb_syn.char_path[70] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02748_));
 sky130_fd_sc_hd__a22o_1 _05691_ (.A1(\top.cb_syn.char_path[38] ),
    .A2(net529),
    .B1(net310),
    .B2(\top.cb_syn.char_path[102] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02749_));
 sky130_fd_sc_hd__or2_1 _05692_ (.A(_02748_),
    .B(_02749_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02750_));
 sky130_fd_sc_hd__a22o_1 _05693_ (.A1(\top.hTree.node_reg[38] ),
    .A2(net307),
    .B1(_02750_),
    .B2(net469),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02751_));
 sky130_fd_sc_hd__a221o_1 _05694_ (.A1(\top.histogram.sram_out[6] ),
    .A2(net358),
    .B1(net408),
    .B2(\top.hTree.node_reg[6] ),
    .C1(_02751_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02752_));
 sky130_fd_sc_hd__a22o_1 _05695_ (.A1(net1392),
    .A2(net170),
    .B1(_02752_),
    .B2(net209),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02344_));
 sky130_fd_sc_hd__a22o_1 _05696_ (.A1(\top.cb_syn.char_path[5] ),
    .A2(net549),
    .B1(net541),
    .B2(\top.cb_syn.char_path[69] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02753_));
 sky130_fd_sc_hd__a22o_1 _05697_ (.A1(\top.cb_syn.char_path[37] ),
    .A2(net529),
    .B1(net310),
    .B2(\top.cb_syn.char_path[101] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02754_));
 sky130_fd_sc_hd__o21a_1 _05698_ (.A1(_02753_),
    .A2(_02754_),
    .B1(net468),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02755_));
 sky130_fd_sc_hd__a22o_1 _05699_ (.A1(\top.histogram.sram_out[5] ),
    .A2(net357),
    .B1(net409),
    .B2(\top.hTree.node_reg[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02756_));
 sky130_fd_sc_hd__a211o_1 _05700_ (.A1(\top.hTree.node_reg[37] ),
    .A2(net307),
    .B1(_02755_),
    .C1(_02756_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02757_));
 sky130_fd_sc_hd__a22o_1 _05701_ (.A1(net1285),
    .A2(net170),
    .B1(_02757_),
    .B2(net209),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02343_));
 sky130_fd_sc_hd__a22o_1 _05702_ (.A1(\top.cb_syn.char_path[4] ),
    .A2(net549),
    .B1(net541),
    .B2(\top.cb_syn.char_path[68] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02758_));
 sky130_fd_sc_hd__a22o_1 _05703_ (.A1(\top.cb_syn.char_path[36] ),
    .A2(net529),
    .B1(net310),
    .B2(\top.cb_syn.char_path[100] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02759_));
 sky130_fd_sc_hd__or2_1 _05704_ (.A(_02758_),
    .B(_02759_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02760_));
 sky130_fd_sc_hd__a22o_1 _05705_ (.A1(\top.hTree.node_reg[36] ),
    .A2(net307),
    .B1(_02760_),
    .B2(net469),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02761_));
 sky130_fd_sc_hd__a221o_1 _05706_ (.A1(\top.histogram.sram_out[4] ),
    .A2(net357),
    .B1(net408),
    .B2(\top.hTree.node_reg[4] ),
    .C1(_02761_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02762_));
 sky130_fd_sc_hd__a22o_1 _05707_ (.A1(net1290),
    .A2(net170),
    .B1(_02762_),
    .B2(net212),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02342_));
 sky130_fd_sc_hd__a22o_1 _05708_ (.A1(\top.cb_syn.char_path[3] ),
    .A2(net548),
    .B1(net539),
    .B2(\top.cb_syn.char_path[67] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02763_));
 sky130_fd_sc_hd__a22o_1 _05709_ (.A1(\top.cb_syn.char_path[35] ),
    .A2(net529),
    .B1(net310),
    .B2(\top.cb_syn.char_path[99] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02764_));
 sky130_fd_sc_hd__or2_1 _05710_ (.A(_02763_),
    .B(_02764_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02765_));
 sky130_fd_sc_hd__a22o_1 _05711_ (.A1(\top.hTree.node_reg[35] ),
    .A2(net307),
    .B1(_02765_),
    .B2(net469),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02766_));
 sky130_fd_sc_hd__a221o_1 _05712_ (.A1(\top.histogram.sram_out[3] ),
    .A2(net357),
    .B1(net408),
    .B2(\top.hTree.node_reg[3] ),
    .C1(_02766_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02767_));
 sky130_fd_sc_hd__a22o_1 _05713_ (.A1(net1248),
    .A2(net170),
    .B1(_02767_),
    .B2(net209),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02341_));
 sky130_fd_sc_hd__a22o_1 _05714_ (.A1(\top.cb_syn.char_path[2] ),
    .A2(net548),
    .B1(net539),
    .B2(\top.cb_syn.char_path[66] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02768_));
 sky130_fd_sc_hd__a22o_1 _05715_ (.A1(\top.cb_syn.char_path[34] ),
    .A2(net530),
    .B1(net311),
    .B2(\top.cb_syn.char_path[98] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02769_));
 sky130_fd_sc_hd__or2_1 _05716_ (.A(_02768_),
    .B(_02769_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02770_));
 sky130_fd_sc_hd__a22o_1 _05717_ (.A1(\top.hTree.node_reg[34] ),
    .A2(net307),
    .B1(_02770_),
    .B2(net469),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02771_));
 sky130_fd_sc_hd__a221o_1 _05718_ (.A1(\top.histogram.sram_out[2] ),
    .A2(net357),
    .B1(net408),
    .B2(\top.hTree.node_reg[2] ),
    .C1(_02771_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02772_));
 sky130_fd_sc_hd__a22o_1 _05719_ (.A1(net1314),
    .A2(net170),
    .B1(_02772_),
    .B2(net209),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02340_));
 sky130_fd_sc_hd__a22o_1 _05720_ (.A1(\top.cb_syn.char_path[1] ),
    .A2(net548),
    .B1(net539),
    .B2(\top.cb_syn.char_path[65] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02773_));
 sky130_fd_sc_hd__a22o_1 _05721_ (.A1(\top.cb_syn.char_path[33] ),
    .A2(net530),
    .B1(net311),
    .B2(\top.cb_syn.char_path[97] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02774_));
 sky130_fd_sc_hd__o21a_1 _05722_ (.A1(_02773_),
    .A2(_02774_),
    .B1(net467),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02775_));
 sky130_fd_sc_hd__a22o_1 _05723_ (.A1(\top.histogram.sram_out[1] ),
    .A2(net357),
    .B1(net408),
    .B2(\top.hTree.node_reg[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02776_));
 sky130_fd_sc_hd__a211o_1 _05724_ (.A1(\top.hTree.node_reg[33] ),
    .A2(net307),
    .B1(_02775_),
    .C1(_02776_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02777_));
 sky130_fd_sc_hd__a22o_1 _05725_ (.A1(net1274),
    .A2(net170),
    .B1(_02777_),
    .B2(net209),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02339_));
 sky130_fd_sc_hd__a22o_1 _05726_ (.A1(\top.cb_syn.char_path[0] ),
    .A2(net546),
    .B1(net538),
    .B2(\top.cb_syn.char_path[64] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02778_));
 sky130_fd_sc_hd__a22o_1 _05727_ (.A1(\top.cb_syn.char_path[32] ),
    .A2(net528),
    .B1(net309),
    .B2(\top.cb_syn.char_path[96] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02779_));
 sky130_fd_sc_hd__or2_2 _05728_ (.A(_02778_),
    .B(_02779_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02780_));
 sky130_fd_sc_hd__a22o_1 _05729_ (.A1(\top.hTree.node_reg[32] ),
    .A2(net308),
    .B1(_02780_),
    .B2(net469),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02781_));
 sky130_fd_sc_hd__a221o_1 _05730_ (.A1(\top.histogram.sram_out[0] ),
    .A2(net357),
    .B1(net408),
    .B2(\top.hTree.node_reg[0] ),
    .C1(_02781_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02782_));
 sky130_fd_sc_hd__a22o_1 _05731_ (.A1(net1473),
    .A2(net170),
    .B1(_02782_),
    .B2(net209),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02338_));
 sky130_fd_sc_hd__mux2_1 _05732_ (.A0(\top.TRN_char_index[6] ),
    .A1(net35),
    .S(net714),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02337_));
 sky130_fd_sc_hd__mux2_1 _05733_ (.A0(\top.TRN_char_index[5] ),
    .A1(net43),
    .S(net715),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02336_));
 sky130_fd_sc_hd__mux2_1 _05734_ (.A0(\top.TRN_char_index[4] ),
    .A1(net42),
    .S(net715),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02335_));
 sky130_fd_sc_hd__mux2_1 _05735_ (.A0(\top.TRN_char_index[3] ),
    .A1(net41),
    .S(net715),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02334_));
 sky130_fd_sc_hd__mux2_1 _05736_ (.A0(net445),
    .A1(net40),
    .S(net715),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02333_));
 sky130_fd_sc_hd__mux2_1 _05737_ (.A0(\top.TRN_char_index[1] ),
    .A1(net39),
    .S(net715),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02332_));
 sky130_fd_sc_hd__mux2_1 _05738_ (.A0(\top.TRN_char_index[0] ),
    .A1(net38),
    .S(net715),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02331_));
 sky130_fd_sc_hd__or2_1 _05739_ (.A(\top.findLeastValue.histo_index[8] ),
    .B(_02575_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02783_));
 sky130_fd_sc_hd__or2_1 _05740_ (.A(\top.findLeastValue.alternator_timer[1] ),
    .B(\top.findLeastValue.alternator_timer[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02784_));
 sky130_fd_sc_hd__a211o_1 _05741_ (.A1(\top.findLeastValue.alternator_timer[2] ),
    .A2(_02784_),
    .B1(_02783_),
    .C1(\top.findLeastValue.alternator_timer[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02785_));
 sky130_fd_sc_hd__nor2_1 _05742_ (.A(\top.findLeastValue.histo_index[8] ),
    .B(\top.findLeastValue.histo_index[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02786_));
 sky130_fd_sc_hd__or2_2 _05743_ (.A(\top.findLeastValue.histo_index[8] ),
    .B(\top.findLeastValue.histo_index[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02787_));
 sky130_fd_sc_hd__o21ai_1 _05744_ (.A1(\top.findLeastValue.alternator_timer[3] ),
    .A2(\top.findLeastValue.alternator_timer[2] ),
    .B1(net406),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02788_));
 sky130_fd_sc_hd__nand2_1 _05745_ (.A(_02783_),
    .B(_02788_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02789_));
 sky130_fd_sc_hd__o21a_1 _05746_ (.A1(\top.findLeastValue.alternator_timer[2] ),
    .A2(_02784_),
    .B1(\top.findLeastValue.alternator_timer[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02790_));
 sky130_fd_sc_hd__o21a_1 _05747_ (.A1(_02789_),
    .A2(_02790_),
    .B1(_02785_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02791_));
 sky130_fd_sc_hd__o211a_1 _05748_ (.A1(\top.findLeastValue.histo_index[7] ),
    .A2(_02789_),
    .B1(_02791_),
    .C1(_02500_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02792_));
 sky130_fd_sc_hd__o21ai_2 _05749_ (.A1(\top.findLeastValue.startup ),
    .A2(_02792_),
    .B1(net457),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02793_));
 sky130_fd_sc_hd__nor2_1 _05750_ (.A(_02783_),
    .B(_02793_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02794_));
 sky130_fd_sc_hd__nor2_1 _05751_ (.A(net444),
    .B(_02562_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02795_));
 sky130_fd_sc_hd__or2_1 _05752_ (.A(net442),
    .B(_02793_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02796_));
 sky130_fd_sc_hd__or3b_1 _05753_ (.A(\top.sram_interface.write_counter_FLV[1] ),
    .B(\top.sram_interface.write_counter_FLV[0] ),
    .C_N(\top.sram_interface.write_counter_FLV[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02797_));
 sky130_fd_sc_hd__inv_2 _05754_ (.A(_02797_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02798_));
 sky130_fd_sc_hd__and2_1 _05755_ (.A(_02576_),
    .B(_02798_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02799_));
 sky130_fd_sc_hd__nand2_1 _05756_ (.A(_02576_),
    .B(_02798_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02800_));
 sky130_fd_sc_hd__and3b_1 _05757_ (.A_N(_02794_),
    .B(_02796_),
    .C(_02800_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02801_));
 sky130_fd_sc_hd__and3_1 _05758_ (.A(net543),
    .B(net457),
    .C(_02801_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02802_));
 sky130_fd_sc_hd__a211o_1 _05759_ (.A1(net542),
    .A2(_02799_),
    .B1(_02802_),
    .C1(_02562_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02803_));
 sky130_fd_sc_hd__nor2_1 _05760_ (.A(net544),
    .B(net536),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02804_));
 sky130_fd_sc_hd__a221o_2 _05761_ (.A1(net442),
    .A2(net536),
    .B1(_02564_),
    .B2(_02804_),
    .C1(_02803_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02805_));
 sky130_fd_sc_hd__nor2_2 _05762_ (.A(_02564_),
    .B(net162),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02806_));
 sky130_fd_sc_hd__a22o_1 _05763_ (.A1(net1802),
    .A2(net163),
    .B1(net147),
    .B2(\top.WB.CPU_DAT_O[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02330_));
 sky130_fd_sc_hd__a22o_1 _05764_ (.A1(\top.compVal[44] ),
    .A2(net163),
    .B1(_02806_),
    .B2(\top.WB.CPU_DAT_O[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02329_));
 sky130_fd_sc_hd__a22o_1 _05765_ (.A1(\top.compVal[43] ),
    .A2(net162),
    .B1(_02806_),
    .B2(\top.WB.CPU_DAT_O[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02328_));
 sky130_fd_sc_hd__a22o_1 _05766_ (.A1(\top.compVal[42] ),
    .A2(net163),
    .B1(net147),
    .B2(\top.WB.CPU_DAT_O[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02327_));
 sky130_fd_sc_hd__a22o_1 _05767_ (.A1(\top.compVal[41] ),
    .A2(net163),
    .B1(_02806_),
    .B2(\top.WB.CPU_DAT_O[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02326_));
 sky130_fd_sc_hd__a22o_1 _05768_ (.A1(\top.compVal[40] ),
    .A2(net163),
    .B1(_02806_),
    .B2(\top.WB.CPU_DAT_O[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02325_));
 sky130_fd_sc_hd__a22o_1 _05769_ (.A1(\top.compVal[39] ),
    .A2(net162),
    .B1(net147),
    .B2(\top.WB.CPU_DAT_O[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02324_));
 sky130_fd_sc_hd__a22o_1 _05770_ (.A1(\top.compVal[38] ),
    .A2(net162),
    .B1(net147),
    .B2(\top.WB.CPU_DAT_O[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02323_));
 sky130_fd_sc_hd__a22o_1 _05771_ (.A1(\top.compVal[37] ),
    .A2(net162),
    .B1(net147),
    .B2(\top.WB.CPU_DAT_O[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02322_));
 sky130_fd_sc_hd__a22o_1 _05772_ (.A1(\top.compVal[36] ),
    .A2(net162),
    .B1(net147),
    .B2(\top.WB.CPU_DAT_O[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02321_));
 sky130_fd_sc_hd__a22o_1 _05773_ (.A1(\top.compVal[35] ),
    .A2(net162),
    .B1(net147),
    .B2(\top.WB.CPU_DAT_O[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02320_));
 sky130_fd_sc_hd__a22o_1 _05774_ (.A1(\top.compVal[34] ),
    .A2(net162),
    .B1(net147),
    .B2(\top.WB.CPU_DAT_O[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02319_));
 sky130_fd_sc_hd__a22o_1 _05775_ (.A1(\top.compVal[33] ),
    .A2(net162),
    .B1(net147),
    .B2(\top.WB.CPU_DAT_O[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02318_));
 sky130_fd_sc_hd__a22o_1 _05776_ (.A1(\top.compVal[32] ),
    .A2(net162),
    .B1(net147),
    .B2(\top.WB.CPU_DAT_O[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02317_));
 sky130_fd_sc_hd__and2_1 _05777_ (.A(net423),
    .B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02807_));
 sky130_fd_sc_hd__and3_1 _05778_ (.A(net423),
    .B(net452),
    .C(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02808_));
 sky130_fd_sc_hd__or4bb_1 _05779_ (.A(net513),
    .B(\top.translation.totalEn ),
    .C_N(_02808_),
    .D_N(\top.TRN_sram_complete ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02809_));
 sky130_fd_sc_hd__or2_2 _05780_ (.A(net506),
    .B(net508),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02810_));
 sky130_fd_sc_hd__nor2_1 _05781_ (.A(net505),
    .B(net402),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02811_));
 sky130_fd_sc_hd__or4_2 _05782_ (.A(\top.translation.index[4] ),
    .B(net502),
    .C(net504),
    .D(net402),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02812_));
 sky130_fd_sc_hd__and3b_1 _05783_ (.A_N(_02812_),
    .B(_02546_),
    .C(_02545_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02813_));
 sky130_fd_sc_hd__or3_1 _05784_ (.A(\top.translation.index[6] ),
    .B(\top.translation.index[5] ),
    .C(_02812_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02814_));
 sky130_fd_sc_hd__nor2_1 _05785_ (.A(_02809_),
    .B(_02814_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02815_));
 sky130_fd_sc_hd__mux2_1 _05786_ (.A0(_02815_),
    .A1(_02809_),
    .S(net1635),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02316_));
 sky130_fd_sc_hd__and2b_1 _05787_ (.A_N(\top.sram_interface.zero_cnt[2] ),
    .B(\top.sram_interface.zero_cnt[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02816_));
 sky130_fd_sc_hd__and2_1 _05788_ (.A(net456),
    .B(\top.sram_interface.word_cnt[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02817_));
 sky130_fd_sc_hd__and3_1 _05789_ (.A(\top.sram_interface.zero_cnt[0] ),
    .B(net456),
    .C(\top.sram_interface.word_cnt[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02818_));
 sky130_fd_sc_hd__nand2b_1 _05790_ (.A_N(_02816_),
    .B(_02818_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02819_));
 sky130_fd_sc_hd__and3_1 _05791_ (.A(\top.sram_interface.zero_cnt[2] ),
    .B(\top.sram_interface.zero_cnt[1] ),
    .C(_02818_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02820_));
 sky130_fd_sc_hd__and2b_1 _05792_ (.A_N(_02820_),
    .B(net1390),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02297_));
 sky130_fd_sc_hd__o21ba_1 _05793_ (.A1(net1489),
    .A2(_02818_),
    .B1_N(_02820_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02296_));
 sky130_fd_sc_hd__o21a_1 _05794_ (.A1(net1428),
    .A2(_02817_),
    .B1(_02819_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02295_));
 sky130_fd_sc_hd__o21a_1 _05795_ (.A1(net1531),
    .A2(net454),
    .B1(_02594_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02294_));
 sky130_fd_sc_hd__o21ai_1 _05796_ (.A1(net542),
    .A2(_02577_),
    .B1(_02800_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02821_));
 sky130_fd_sc_hd__nand2_1 _05797_ (.A(net444),
    .B(net527),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02822_));
 sky130_fd_sc_hd__o311a_1 _05798_ (.A1(net542),
    .A2(net533),
    .A3(net527),
    .B1(_02821_),
    .C1(_02822_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02823_));
 sky130_fd_sc_hd__nand2_1 _05799_ (.A(net455),
    .B(_02823_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02824_));
 sky130_fd_sc_hd__o211a_1 _05800_ (.A1(net533),
    .A2(net527),
    .B1(_02823_),
    .C1(net455),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02825_));
 sky130_fd_sc_hd__nand2_1 _05801_ (.A(\top.sram_interface.write_counter_FLV[1] ),
    .B(\top.sram_interface.write_counter_FLV[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02826_));
 sky130_fd_sc_hd__xnor2_1 _05802_ (.A(\top.sram_interface.write_counter_FLV[2] ),
    .B(_02826_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02827_));
 sky130_fd_sc_hd__a22o_1 _05803_ (.A1(net1631),
    .A2(_02824_),
    .B1(_02825_),
    .B2(_02827_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02293_));
 sky130_fd_sc_hd__nand3_1 _05804_ (.A(\top.sram_interface.write_counter_FLV[0] ),
    .B(net455),
    .C(_02823_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02828_));
 sky130_fd_sc_hd__xnor2_1 _05805_ (.A(net1281),
    .B(_02828_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02292_));
 sky130_fd_sc_hd__o21a_1 _05806_ (.A1(net1633),
    .A2(_02825_),
    .B1(_02828_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02291_));
 sky130_fd_sc_hd__or4_1 _05807_ (.A(\top.findLeastValue.least1[3] ),
    .B(\top.findLeastValue.least1[2] ),
    .C(\top.findLeastValue.least1[1] ),
    .D(\top.findLeastValue.least1[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02829_));
 sky130_fd_sc_hd__or4_1 _05808_ (.A(_02523_),
    .B(\top.findLeastValue.least1[6] ),
    .C(\top.findLeastValue.least1[5] ),
    .D(\top.findLeastValue.least1[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02830_));
 sky130_fd_sc_hd__nor2_1 _05809_ (.A(_02829_),
    .B(_02830_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02831_));
 sky130_fd_sc_hd__nand2_1 _05810_ (.A(\top.findLeastValue.least1[8] ),
    .B(_02831_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02832_));
 sky130_fd_sc_hd__or4_1 _05811_ (.A(\top.findLeastValue.least2[3] ),
    .B(\top.findLeastValue.least2[2] ),
    .C(\top.findLeastValue.least2[1] ),
    .D(\top.findLeastValue.least2[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02833_));
 sky130_fd_sc_hd__or4b_1 _05812_ (.A(\top.findLeastValue.least2[6] ),
    .B(\top.findLeastValue.least2[5] ),
    .C(\top.findLeastValue.least2[4] ),
    .D_N(\top.findLeastValue.least2[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02834_));
 sky130_fd_sc_hd__nor2_1 _05813_ (.A(_02833_),
    .B(_02834_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02835_));
 sky130_fd_sc_hd__nand2_1 _05814_ (.A(\top.findLeastValue.least2[8] ),
    .B(_02835_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02836_));
 sky130_fd_sc_hd__or2_2 _05815_ (.A(_02832_),
    .B(_02836_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02837_));
 sky130_fd_sc_hd__or3b_1 _05816_ (.A(\top.hTree.write_HT_fin ),
    .B(net417),
    .C_N(_02837_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02838_));
 sky130_fd_sc_hd__nor2_1 _05817_ (.A(net442),
    .B(net431),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02839_));
 sky130_fd_sc_hd__or3_1 _05818_ (.A(net442),
    .B(net431),
    .C(_02838_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02840_));
 sky130_fd_sc_hd__nor3_1 _05819_ (.A(net442),
    .B(\top.sram_interface.counter_HTREE[3] ),
    .C(\top.sram_interface.counter_HTREE[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02841_));
 sky130_fd_sc_hd__and3b_1 _05820_ (.A_N(\top.sram_interface.counter_HTREE[0] ),
    .B(_02841_),
    .C(\top.sram_interface.counter_HTREE[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02842_));
 sky130_fd_sc_hd__or3b_1 _05821_ (.A(\top.findLeastValue.least2[8] ),
    .B(\top.findLeastValue.least1[8] ),
    .C_N(_02842_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02843_));
 sky130_fd_sc_hd__nand2_1 _05822_ (.A(_02840_),
    .B(_02843_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02844_));
 sky130_fd_sc_hd__inv_2 _05823_ (.A(_02844_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02845_));
 sky130_fd_sc_hd__nor2_1 _05824_ (.A(\top.hTree.state[6] ),
    .B(\top.hTree.state[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02846_));
 sky130_fd_sc_hd__nand2b_1 _05825_ (.A_N(_02846_),
    .B(_02842_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02847_));
 sky130_fd_sc_hd__or2_1 _05826_ (.A(\top.sram_interface.counter_HTREE[1] ),
    .B(\top.sram_interface.counter_HTREE[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02848_));
 sky130_fd_sc_hd__or3b_1 _05827_ (.A(_02848_),
    .B(\top.sram_interface.counter_HTREE[3] ),
    .C_N(\top.sram_interface.counter_HTREE[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02849_));
 sky130_fd_sc_hd__nor2_1 _05828_ (.A(\top.hTree.state[7] ),
    .B(\top.hTree.state[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02850_));
 sky130_fd_sc_hd__or2_2 _05829_ (.A(\top.hTree.state[7] ),
    .B(\top.hTree.state[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02851_));
 sky130_fd_sc_hd__or3_1 _05830_ (.A(net443),
    .B(_02849_),
    .C(net401),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02852_));
 sky130_fd_sc_hd__nor2_1 _05831_ (.A(_02514_),
    .B(_02522_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02853_));
 sky130_fd_sc_hd__and2_1 _05832_ (.A(\top.sram_interface.counter_HTREE[1] ),
    .B(\top.sram_interface.counter_HTREE[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02854_));
 sky130_fd_sc_hd__nand2_1 _05833_ (.A(\top.sram_interface.counter_HTREE[1] ),
    .B(\top.sram_interface.counter_HTREE[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02855_));
 sky130_fd_sc_hd__and4_1 _05834_ (.A(\top.hTree.state[2] ),
    .B(_02841_),
    .C(_02853_),
    .D(_02854_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02856_));
 sky130_fd_sc_hd__and4bb_1 _05835_ (.A_N(\top.WorR ),
    .B_N(_02856_),
    .C(net544),
    .D(_02847_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02857_));
 sky130_fd_sc_hd__and4_1 _05836_ (.A(net448),
    .B(_02845_),
    .C(_02852_),
    .D(_02857_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02858_));
 sky130_fd_sc_hd__or4_1 _05837_ (.A(\top.WorR ),
    .B(_02553_),
    .C(_02844_),
    .D(_02847_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02859_));
 sky130_fd_sc_hd__inv_2 _05838_ (.A(_02859_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02860_));
 sky130_fd_sc_hd__or4_2 _05839_ (.A(\top.sram_interface.word_cnt[12] ),
    .B(net533),
    .C(net536),
    .D(\top.sram_interface.word_cnt[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02861_));
 sky130_fd_sc_hd__o31a_1 _05840_ (.A1(net526),
    .A2(net536),
    .A3(\top.sram_interface.word_cnt[13] ),
    .B1(net446),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02862_));
 sky130_fd_sc_hd__o21ai_1 _05841_ (.A1(net544),
    .A2(_02861_),
    .B1(net448),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02863_));
 sky130_fd_sc_hd__and4b_1 _05842_ (.A_N(_02849_),
    .B(net440),
    .C(\top.hTree.state[8] ),
    .D(_02853_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02864_));
 sky130_fd_sc_hd__and3_1 _05843_ (.A(_02832_),
    .B(_02836_),
    .C(_02864_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02865_));
 sky130_fd_sc_hd__and3_1 _05844_ (.A(net448),
    .B(net544),
    .C(_02865_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02866_));
 sky130_fd_sc_hd__or4_2 _05845_ (.A(_02858_),
    .B(_02860_),
    .C(_02863_),
    .D(_02866_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02867_));
 sky130_fd_sc_hd__nand2_1 _05846_ (.A(\top.sram_interface.counter_HTREE[2] ),
    .B(_02854_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02868_));
 sky130_fd_sc_hd__a21o_1 _05847_ (.A1(_02861_),
    .A2(_02868_),
    .B1(_02867_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02869_));
 sky130_fd_sc_hd__and2b_1 _05848_ (.A_N(_02867_),
    .B(_02861_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02870_));
 sky130_fd_sc_hd__nor2_1 _05849_ (.A(\top.sram_interface.counter_HTREE[3] ),
    .B(_02868_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02871_));
 sky130_fd_sc_hd__a22o_1 _05850_ (.A1(net1761),
    .A2(_02869_),
    .B1(_02870_),
    .B2(_02871_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02290_));
 sky130_fd_sc_hd__nor2_1 _05851_ (.A(_02855_),
    .B(_02867_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02872_));
 sky130_fd_sc_hd__o21a_1 _05852_ (.A1(net1640),
    .A2(_02872_),
    .B1(_02869_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02289_));
 sky130_fd_sc_hd__a32o_1 _05853_ (.A1(_02848_),
    .A2(_02855_),
    .A3(_02870_),
    .B1(_02867_),
    .B2(net1690),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02288_));
 sky130_fd_sc_hd__mux2_1 _05854_ (.A0(_02870_),
    .A1(_02867_),
    .S(\top.sram_interface.counter_HTREE[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02287_));
 sky130_fd_sc_hd__or4_1 _05855_ (.A(\top.sram_interface.init_counter[15] ),
    .B(\top.sram_interface.init_counter[14] ),
    .C(\top.sram_interface.init_counter[13] ),
    .D(\top.sram_interface.init_counter[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02873_));
 sky130_fd_sc_hd__or4_1 _05856_ (.A(\top.sram_interface.init_counter[19] ),
    .B(\top.sram_interface.init_counter[18] ),
    .C(\top.sram_interface.init_counter[17] ),
    .D(\top.sram_interface.init_counter[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02874_));
 sky130_fd_sc_hd__or4_1 _05857_ (.A(\top.sram_interface.init_counter[23] ),
    .B(\top.sram_interface.init_counter[22] ),
    .C(\top.sram_interface.init_counter[21] ),
    .D(\top.sram_interface.init_counter[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02875_));
 sky130_fd_sc_hd__or3_1 _05858_ (.A(_02873_),
    .B(_02874_),
    .C(_02875_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02876_));
 sky130_fd_sc_hd__nor2_1 _05859_ (.A(\top.sram_interface.init_counter[11] ),
    .B(_02876_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02877_));
 sky130_fd_sc_hd__and3_1 _05860_ (.A(net439),
    .B(\top.WB.prev_BUSY_O ),
    .C(_02877_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02878_));
 sky130_fd_sc_hd__o31a_1 _05861_ (.A1(_02417_),
    .A2(_02447_),
    .A3(_02878_),
    .B1(net481),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02286_));
 sky130_fd_sc_hd__or3_1 _05862_ (.A(_02553_),
    .B(_02562_),
    .C(_02801_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02879_));
 sky130_fd_sc_hd__and3_1 _05863_ (.A(net542),
    .B(net456),
    .C(_02799_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02880_));
 sky130_fd_sc_hd__a21o_1 _05864_ (.A1(net1476),
    .A2(_02879_),
    .B1(_02880_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02285_));
 sky130_fd_sc_hd__o22a_1 _05865_ (.A1(net448),
    .A2(_02562_),
    .B1(net411),
    .B2(\top.hTree.write_HT_fin ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02284_));
 sky130_fd_sc_hd__and3_1 _05866_ (.A(net439),
    .B(net453),
    .C(\top.histogram.state[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02881_));
 sky130_fd_sc_hd__mux2_1 _05867_ (.A0(net1526),
    .A1(\top.WB.CPU_DAT_O[31] ),
    .S(net353),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02283_));
 sky130_fd_sc_hd__mux2_1 _05868_ (.A0(net1646),
    .A1(\top.WB.CPU_DAT_O[30] ),
    .S(net353),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02282_));
 sky130_fd_sc_hd__mux2_1 _05869_ (.A0(net1529),
    .A1(\top.WB.CPU_DAT_O[29] ),
    .S(net353),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02281_));
 sky130_fd_sc_hd__mux2_1 _05870_ (.A0(net1524),
    .A1(\top.WB.CPU_DAT_O[28] ),
    .S(net353),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02280_));
 sky130_fd_sc_hd__mux2_1 _05871_ (.A0(net1774),
    .A1(\top.WB.CPU_DAT_O[27] ),
    .S(net350),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02279_));
 sky130_fd_sc_hd__mux2_1 _05872_ (.A0(net1509),
    .A1(\top.WB.CPU_DAT_O[26] ),
    .S(net350),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02278_));
 sky130_fd_sc_hd__mux2_1 _05873_ (.A0(net1481),
    .A1(\top.WB.CPU_DAT_O[25] ),
    .S(net350),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02277_));
 sky130_fd_sc_hd__mux2_1 _05874_ (.A0(\top.hist_data_o[24] ),
    .A1(\top.WB.CPU_DAT_O[24] ),
    .S(net350),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02276_));
 sky130_fd_sc_hd__mux2_1 _05875_ (.A0(net1388),
    .A1(\top.WB.CPU_DAT_O[23] ),
    .S(net350),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02275_));
 sky130_fd_sc_hd__mux2_1 _05876_ (.A0(net1536),
    .A1(\top.WB.CPU_DAT_O[22] ),
    .S(net350),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02274_));
 sky130_fd_sc_hd__mux2_1 _05877_ (.A0(net1625),
    .A1(\top.WB.CPU_DAT_O[21] ),
    .S(net350),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02273_));
 sky130_fd_sc_hd__mux2_1 _05878_ (.A0(net1760),
    .A1(\top.WB.CPU_DAT_O[20] ),
    .S(net350),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02272_));
 sky130_fd_sc_hd__mux2_1 _05879_ (.A0(net1718),
    .A1(\top.WB.CPU_DAT_O[19] ),
    .S(net350),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02271_));
 sky130_fd_sc_hd__mux2_1 _05880_ (.A0(net1686),
    .A1(\top.WB.CPU_DAT_O[18] ),
    .S(net350),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02270_));
 sky130_fd_sc_hd__mux2_1 _05881_ (.A0(net1663),
    .A1(\top.WB.CPU_DAT_O[17] ),
    .S(net351),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02269_));
 sky130_fd_sc_hd__mux2_1 _05882_ (.A0(net1689),
    .A1(\top.WB.CPU_DAT_O[16] ),
    .S(net351),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02268_));
 sky130_fd_sc_hd__mux2_1 _05883_ (.A0(net1790),
    .A1(\top.WB.CPU_DAT_O[15] ),
    .S(net351),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02267_));
 sky130_fd_sc_hd__mux2_1 _05884_ (.A0(net1606),
    .A1(\top.WB.CPU_DAT_O[14] ),
    .S(net351),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02266_));
 sky130_fd_sc_hd__mux2_1 _05885_ (.A0(net1562),
    .A1(\top.WB.CPU_DAT_O[13] ),
    .S(net351),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02265_));
 sky130_fd_sc_hd__mux2_1 _05886_ (.A0(net1623),
    .A1(\top.WB.CPU_DAT_O[12] ),
    .S(net351),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02264_));
 sky130_fd_sc_hd__mux2_1 _05887_ (.A0(net1534),
    .A1(\top.WB.CPU_DAT_O[11] ),
    .S(net349),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02263_));
 sky130_fd_sc_hd__mux2_1 _05888_ (.A0(net1634),
    .A1(\top.WB.CPU_DAT_O[10] ),
    .S(net349),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02262_));
 sky130_fd_sc_hd__mux2_1 _05889_ (.A0(\top.hist_data_o[9] ),
    .A1(\top.WB.CPU_DAT_O[9] ),
    .S(net352),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02261_));
 sky130_fd_sc_hd__mux2_1 _05890_ (.A0(\top.hist_data_o[8] ),
    .A1(\top.WB.CPU_DAT_O[8] ),
    .S(net352),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02260_));
 sky130_fd_sc_hd__mux2_1 _05891_ (.A0(net1549),
    .A1(\top.WB.CPU_DAT_O[7] ),
    .S(net349),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02259_));
 sky130_fd_sc_hd__mux2_1 _05892_ (.A0(\top.hist_data_o[6] ),
    .A1(\top.WB.CPU_DAT_O[6] ),
    .S(net349),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02258_));
 sky130_fd_sc_hd__mux2_1 _05893_ (.A0(net1528),
    .A1(\top.WB.CPU_DAT_O[5] ),
    .S(net349),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02257_));
 sky130_fd_sc_hd__mux2_1 _05894_ (.A0(\top.hist_data_o[4] ),
    .A1(\top.WB.CPU_DAT_O[4] ),
    .S(net349),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02256_));
 sky130_fd_sc_hd__mux2_1 _05895_ (.A0(net1577),
    .A1(\top.WB.CPU_DAT_O[3] ),
    .S(net349),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02255_));
 sky130_fd_sc_hd__mux2_1 _05896_ (.A0(\top.hist_data_o[2] ),
    .A1(\top.WB.CPU_DAT_O[2] ),
    .S(net349),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02254_));
 sky130_fd_sc_hd__mux2_1 _05897_ (.A0(\top.hist_data_o[1] ),
    .A1(\top.WB.CPU_DAT_O[1] ),
    .S(net349),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02253_));
 sky130_fd_sc_hd__mux2_1 _05898_ (.A0(\top.hist_data_o[0] ),
    .A1(\top.WB.CPU_DAT_O[0] ),
    .S(net349),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02252_));
 sky130_fd_sc_hd__a21o_1 _05899_ (.A1(net461),
    .A2(\top.sram_interface.word_cnt[9] ),
    .B1(net956),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02251_));
 sky130_fd_sc_hd__or4_1 _05900_ (.A(\top.cb_syn.h_element[49] ),
    .B(\top.cb_syn.h_element[48] ),
    .C(\top.cb_syn.h_element[47] ),
    .D(\top.cb_syn.h_element[46] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02882_));
 sky130_fd_sc_hd__or4b_1 _05901_ (.A(\top.cb_syn.h_element[52] ),
    .B(\top.cb_syn.h_element[51] ),
    .C(\top.cb_syn.h_element[50] ),
    .D_N(\top.cb_syn.h_element[53] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02883_));
 sky130_fd_sc_hd__o21ai_1 _05902_ (.A1(_02882_),
    .A2(_02883_),
    .B1(\top.cb_syn.h_element[54] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02884_));
 sky130_fd_sc_hd__or2_1 _05903_ (.A(net489),
    .B(_02538_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02885_));
 sky130_fd_sc_hd__inv_2 _05904_ (.A(_02885_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02886_));
 sky130_fd_sc_hd__nor2_1 _05905_ (.A(_02884_),
    .B(_02885_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02887_));
 sky130_fd_sc_hd__and2b_1 _05906_ (.A_N(\top.cb_syn.end_check ),
    .B(\top.cb_syn.curr_state[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02888_));
 sky130_fd_sc_hd__nor2_1 _05907_ (.A(net488),
    .B(net412),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02889_));
 sky130_fd_sc_hd__or2_1 _05908_ (.A(net488),
    .B(net412),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02890_));
 sky130_fd_sc_hd__nand2_1 _05909_ (.A(net521),
    .B(_02889_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02891_));
 sky130_fd_sc_hd__or4_1 _05910_ (.A(\top.cb_syn.h_element[58] ),
    .B(\top.cb_syn.h_element[57] ),
    .C(\top.cb_syn.h_element[56] ),
    .D(\top.cb_syn.h_element[55] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02892_));
 sky130_fd_sc_hd__or4b_1 _05911_ (.A(\top.cb_syn.h_element[61] ),
    .B(\top.cb_syn.h_element[60] ),
    .C(\top.cb_syn.h_element[59] ),
    .D_N(\top.cb_syn.h_element[62] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02893_));
 sky130_fd_sc_hd__nor2_1 _05912_ (.A(_02892_),
    .B(_02893_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02894_));
 sky130_fd_sc_hd__nor2_1 _05913_ (.A(_02551_),
    .B(_02894_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02895_));
 sky130_fd_sc_hd__and3b_1 _05914_ (.A_N(net489),
    .B(net524),
    .C(_02895_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02896_));
 sky130_fd_sc_hd__o21ai_1 _05915_ (.A1(_02887_),
    .A2(_02896_),
    .B1(_02581_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02897_));
 sky130_fd_sc_hd__and3b_1 _05916_ (.A_N(_02888_),
    .B(_02891_),
    .C(_02897_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02898_));
 sky130_fd_sc_hd__and3_1 _05917_ (.A(net439),
    .B(net543),
    .C(net460),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02899_));
 sky130_fd_sc_hd__nor2_1 _05918_ (.A(net442),
    .B(_02898_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02900_));
 sky130_fd_sc_hd__or2_1 _05919_ (.A(net442),
    .B(_02898_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02901_));
 sky130_fd_sc_hd__and3_1 _05920_ (.A(net542),
    .B(net460),
    .C(_02900_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02902_));
 sky130_fd_sc_hd__a31o_1 _05921_ (.A1(_02553_),
    .A2(net460),
    .A3(_02588_),
    .B1(_02902_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02903_));
 sky130_fd_sc_hd__o21ai_1 _05922_ (.A1(\top.sram_interface.CB_write_counter[0] ),
    .A2(_02587_),
    .B1(_02903_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02904_));
 sky130_fd_sc_hd__nor2_1 _05923_ (.A(\top.sram_interface.CB_write_counter[1] ),
    .B(_02587_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02905_));
 sky130_fd_sc_hd__a32o_1 _05924_ (.A1(\top.sram_interface.CB_write_counter[0] ),
    .A2(_02903_),
    .A3(_02905_),
    .B1(_02904_),
    .B2(\top.sram_interface.CB_write_counter[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02250_));
 sky130_fd_sc_hd__o21a_1 _05925_ (.A1(\top.sram_interface.CB_write_counter[0] ),
    .A2(_02903_),
    .B1(_02904_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02249_));
 sky130_fd_sc_hd__nor2_1 _05926_ (.A(net536),
    .B(net537),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02906_));
 sky130_fd_sc_hd__mux2_1 _05927_ (.A0(net443),
    .A1(_02553_),
    .S(_02906_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02907_));
 sky130_fd_sc_hd__or2_2 _05928_ (.A(_02803_),
    .B(_02907_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02908_));
 sky130_fd_sc_hd__nor2_1 _05929_ (.A(_02906_),
    .B(net158),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02909_));
 sky130_fd_sc_hd__a22o_1 _05930_ (.A1(\top.compVal[31] ),
    .A2(net159),
    .B1(net144),
    .B2(\top.WB.CPU_DAT_O[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02248_));
 sky130_fd_sc_hd__a22o_1 _05931_ (.A1(\top.compVal[30] ),
    .A2(net158),
    .B1(net145),
    .B2(\top.WB.CPU_DAT_O[30] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02247_));
 sky130_fd_sc_hd__a22o_1 _05932_ (.A1(\top.compVal[29] ),
    .A2(net158),
    .B1(net145),
    .B2(\top.WB.CPU_DAT_O[29] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02246_));
 sky130_fd_sc_hd__a22o_1 _05933_ (.A1(\top.compVal[28] ),
    .A2(net159),
    .B1(net144),
    .B2(\top.WB.CPU_DAT_O[28] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02245_));
 sky130_fd_sc_hd__a22o_1 _05934_ (.A1(\top.compVal[27] ),
    .A2(net158),
    .B1(net145),
    .B2(\top.WB.CPU_DAT_O[27] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02244_));
 sky130_fd_sc_hd__a22o_1 _05935_ (.A1(\top.compVal[26] ),
    .A2(net158),
    .B1(net146),
    .B2(\top.WB.CPU_DAT_O[26] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02243_));
 sky130_fd_sc_hd__a22o_1 _05936_ (.A1(\top.compVal[25] ),
    .A2(net158),
    .B1(net146),
    .B2(\top.WB.CPU_DAT_O[25] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02242_));
 sky130_fd_sc_hd__a22o_1 _05937_ (.A1(net1127),
    .A2(net158),
    .B1(net145),
    .B2(\top.WB.CPU_DAT_O[24] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02241_));
 sky130_fd_sc_hd__a22o_1 _05938_ (.A1(\top.compVal[23] ),
    .A2(net159),
    .B1(net145),
    .B2(\top.WB.CPU_DAT_O[23] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02240_));
 sky130_fd_sc_hd__a22o_1 _05939_ (.A1(\top.compVal[22] ),
    .A2(net158),
    .B1(net145),
    .B2(\top.WB.CPU_DAT_O[22] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02239_));
 sky130_fd_sc_hd__a22o_1 _05940_ (.A1(\top.compVal[21] ),
    .A2(net158),
    .B1(net145),
    .B2(\top.WB.CPU_DAT_O[21] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02238_));
 sky130_fd_sc_hd__a22o_1 _05941_ (.A1(\top.compVal[20] ),
    .A2(net159),
    .B1(net145),
    .B2(\top.WB.CPU_DAT_O[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02237_));
 sky130_fd_sc_hd__a22o_1 _05942_ (.A1(\top.compVal[19] ),
    .A2(net159),
    .B1(net145),
    .B2(\top.WB.CPU_DAT_O[19] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02236_));
 sky130_fd_sc_hd__a22o_1 _05943_ (.A1(\top.compVal[18] ),
    .A2(net158),
    .B1(net145),
    .B2(\top.WB.CPU_DAT_O[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02235_));
 sky130_fd_sc_hd__a22o_1 _05944_ (.A1(\top.compVal[17] ),
    .A2(net161),
    .B1(net146),
    .B2(\top.WB.CPU_DAT_O[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02234_));
 sky130_fd_sc_hd__a22o_1 _05945_ (.A1(\top.compVal[16] ),
    .A2(net161),
    .B1(net146),
    .B2(\top.WB.CPU_DAT_O[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02233_));
 sky130_fd_sc_hd__a22o_1 _05946_ (.A1(\top.compVal[15] ),
    .A2(net161),
    .B1(net146),
    .B2(\top.WB.CPU_DAT_O[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02232_));
 sky130_fd_sc_hd__a22o_1 _05947_ (.A1(\top.compVal[14] ),
    .A2(net161),
    .B1(net146),
    .B2(\top.WB.CPU_DAT_O[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02231_));
 sky130_fd_sc_hd__a22o_1 _05948_ (.A1(\top.compVal[13] ),
    .A2(net161),
    .B1(net146),
    .B2(\top.WB.CPU_DAT_O[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02230_));
 sky130_fd_sc_hd__a22o_1 _05949_ (.A1(\top.compVal[12] ),
    .A2(net161),
    .B1(net146),
    .B2(\top.WB.CPU_DAT_O[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02229_));
 sky130_fd_sc_hd__a22o_1 _05950_ (.A1(\top.compVal[11] ),
    .A2(net160),
    .B1(net143),
    .B2(\top.WB.CPU_DAT_O[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02228_));
 sky130_fd_sc_hd__a22o_1 _05951_ (.A1(\top.compVal[10] ),
    .A2(net160),
    .B1(net143),
    .B2(\top.WB.CPU_DAT_O[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02227_));
 sky130_fd_sc_hd__a22o_1 _05952_ (.A1(\top.compVal[9] ),
    .A2(net161),
    .B1(net144),
    .B2(\top.WB.CPU_DAT_O[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02226_));
 sky130_fd_sc_hd__a22o_1 _05953_ (.A1(\top.compVal[8] ),
    .A2(net161),
    .B1(net144),
    .B2(\top.WB.CPU_DAT_O[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02225_));
 sky130_fd_sc_hd__a22o_1 _05954_ (.A1(\top.compVal[7] ),
    .A2(net160),
    .B1(net143),
    .B2(\top.WB.CPU_DAT_O[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02224_));
 sky130_fd_sc_hd__a22o_1 _05955_ (.A1(\top.compVal[6] ),
    .A2(net160),
    .B1(net143),
    .B2(\top.WB.CPU_DAT_O[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02223_));
 sky130_fd_sc_hd__a22o_1 _05956_ (.A1(\top.compVal[5] ),
    .A2(net160),
    .B1(net143),
    .B2(\top.WB.CPU_DAT_O[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02222_));
 sky130_fd_sc_hd__a22o_1 _05957_ (.A1(\top.compVal[4] ),
    .A2(net160),
    .B1(net143),
    .B2(\top.WB.CPU_DAT_O[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02221_));
 sky130_fd_sc_hd__a22o_1 _05958_ (.A1(\top.compVal[3] ),
    .A2(net160),
    .B1(net143),
    .B2(\top.WB.CPU_DAT_O[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02220_));
 sky130_fd_sc_hd__a22o_1 _05959_ (.A1(net1804),
    .A2(net160),
    .B1(net143),
    .B2(\top.WB.CPU_DAT_O[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02219_));
 sky130_fd_sc_hd__a22o_1 _05960_ (.A1(\top.compVal[1] ),
    .A2(net160),
    .B1(net143),
    .B2(\top.WB.CPU_DAT_O[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02218_));
 sky130_fd_sc_hd__a22o_1 _05961_ (.A1(\top.compVal[0] ),
    .A2(net160),
    .B1(net143),
    .B2(\top.WB.CPU_DAT_O[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02217_));
 sky130_fd_sc_hd__and2b_1 _05962_ (.A_N(\top.sram_interface.CB_write_counter[0] ),
    .B(\top.sram_interface.CB_write_counter[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02910_));
 sky130_fd_sc_hd__and4b_1 _05963_ (.A_N(_02910_),
    .B(_02899_),
    .C(_02898_),
    .D(\top.sram_interface.CB_read_counter ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02911_));
 sky130_fd_sc_hd__o21ba_1 _05964_ (.A1(\top.CB_read_complete ),
    .A2(_02911_),
    .B1_N(_02902_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02216_));
 sky130_fd_sc_hd__a21oi_1 _05965_ (.A1(_02899_),
    .A2(_02910_),
    .B1(\top.CB_write_complete ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02912_));
 sky130_fd_sc_hd__nor2_1 _05966_ (.A(_02902_),
    .B(_02912_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02215_));
 sky130_fd_sc_hd__and3b_1 _05967_ (.A_N(\top.sram_interface.TRN_counter[2] ),
    .B(\top.sram_interface.TRN_counter[1] ),
    .C(\top.sram_interface.TRN_counter[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02913_));
 sky130_fd_sc_hd__nand2_1 _05968_ (.A(net452),
    .B(net536),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02914_));
 sky130_fd_sc_hd__nand3_1 _05969_ (.A(net452),
    .B(net536),
    .C(_02913_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02915_));
 sky130_fd_sc_hd__mux2_1 _05970_ (.A0(\top.WB.CPU_DAT_O[31] ),
    .A1(net1399),
    .S(net346),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02214_));
 sky130_fd_sc_hd__mux2_1 _05971_ (.A0(\top.WB.CPU_DAT_O[30] ),
    .A1(net1243),
    .S(net346),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02213_));
 sky130_fd_sc_hd__mux2_1 _05972_ (.A0(\top.WB.CPU_DAT_O[29] ),
    .A1(net1400),
    .S(net345),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02212_));
 sky130_fd_sc_hd__mux2_1 _05973_ (.A0(\top.WB.CPU_DAT_O[28] ),
    .A1(net1375),
    .S(net346),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02211_));
 sky130_fd_sc_hd__mux2_1 _05974_ (.A0(\top.WB.CPU_DAT_O[27] ),
    .A1(net1185),
    .S(net345),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02210_));
 sky130_fd_sc_hd__mux2_1 _05975_ (.A0(\top.WB.CPU_DAT_O[26] ),
    .A1(net1283),
    .S(net345),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02209_));
 sky130_fd_sc_hd__mux2_1 _05976_ (.A0(\top.WB.CPU_DAT_O[25] ),
    .A1(net1172),
    .S(net345),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02208_));
 sky130_fd_sc_hd__mux2_1 _05977_ (.A0(\top.WB.CPU_DAT_O[24] ),
    .A1(net1154),
    .S(net345),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02207_));
 sky130_fd_sc_hd__mux2_1 _05978_ (.A0(\top.WB.CPU_DAT_O[23] ),
    .A1(net1227),
    .S(net345),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02206_));
 sky130_fd_sc_hd__mux2_1 _05979_ (.A0(\top.WB.CPU_DAT_O[22] ),
    .A1(net1296),
    .S(net345),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02205_));
 sky130_fd_sc_hd__mux2_1 _05980_ (.A0(\top.WB.CPU_DAT_O[21] ),
    .A1(net1051),
    .S(net345),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02204_));
 sky130_fd_sc_hd__mux2_1 _05981_ (.A0(\top.WB.CPU_DAT_O[20] ),
    .A1(net1219),
    .S(net345),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02203_));
 sky130_fd_sc_hd__mux2_1 _05982_ (.A0(\top.WB.CPU_DAT_O[19] ),
    .A1(net1189),
    .S(net346),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02202_));
 sky130_fd_sc_hd__mux2_1 _05983_ (.A0(\top.WB.CPU_DAT_O[18] ),
    .A1(net1117),
    .S(net346),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02201_));
 sky130_fd_sc_hd__mux2_1 _05984_ (.A0(\top.WB.CPU_DAT_O[17] ),
    .A1(net1391),
    .S(net346),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02200_));
 sky130_fd_sc_hd__mux2_1 _05985_ (.A0(\top.WB.CPU_DAT_O[16] ),
    .A1(net1299),
    .S(net345),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02199_));
 sky130_fd_sc_hd__mux2_1 _05986_ (.A0(\top.WB.CPU_DAT_O[15] ),
    .A1(net1236),
    .S(net347),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02198_));
 sky130_fd_sc_hd__mux2_1 _05987_ (.A0(\top.WB.CPU_DAT_O[14] ),
    .A1(net1256),
    .S(net347),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02197_));
 sky130_fd_sc_hd__mux2_1 _05988_ (.A0(\top.WB.CPU_DAT_O[13] ),
    .A1(net1441),
    .S(net348),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02196_));
 sky130_fd_sc_hd__mux2_1 _05989_ (.A0(\top.WB.CPU_DAT_O[12] ),
    .A1(net1208),
    .S(net348),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02195_));
 sky130_fd_sc_hd__mux2_1 _05990_ (.A0(\top.WB.CPU_DAT_O[11] ),
    .A1(net1150),
    .S(net348),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02194_));
 sky130_fd_sc_hd__mux2_1 _05991_ (.A0(\top.WB.CPU_DAT_O[10] ),
    .A1(net1059),
    .S(net348),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02193_));
 sky130_fd_sc_hd__mux2_1 _05992_ (.A0(\top.WB.CPU_DAT_O[9] ),
    .A1(net1332),
    .S(net347),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02192_));
 sky130_fd_sc_hd__mux2_1 _05993_ (.A0(\top.WB.CPU_DAT_O[8] ),
    .A1(net1201),
    .S(net347),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02191_));
 sky130_fd_sc_hd__mux2_1 _05994_ (.A0(\top.WB.CPU_DAT_O[7] ),
    .A1(net1076),
    .S(net347),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02190_));
 sky130_fd_sc_hd__mux2_1 _05995_ (.A0(\top.WB.CPU_DAT_O[6] ),
    .A1(net1142),
    .S(net347),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02189_));
 sky130_fd_sc_hd__mux2_1 _05996_ (.A0(\top.WB.CPU_DAT_O[5] ),
    .A1(net1052),
    .S(net347),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02188_));
 sky130_fd_sc_hd__mux2_1 _05997_ (.A0(\top.WB.CPU_DAT_O[4] ),
    .A1(net1166),
    .S(net348),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02187_));
 sky130_fd_sc_hd__mux2_1 _05998_ (.A0(\top.WB.CPU_DAT_O[3] ),
    .A1(net1412),
    .S(net347),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02186_));
 sky130_fd_sc_hd__mux2_1 _05999_ (.A0(\top.WB.CPU_DAT_O[2] ),
    .A1(net1138),
    .S(net347),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02185_));
 sky130_fd_sc_hd__mux2_1 _06000_ (.A0(\top.WB.CPU_DAT_O[1] ),
    .A1(net1339),
    .S(net347),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02184_));
 sky130_fd_sc_hd__mux2_1 _06001_ (.A0(\top.WB.CPU_DAT_O[0] ),
    .A1(net1343),
    .S(net348),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02183_));
 sky130_fd_sc_hd__nand2_1 _06002_ (.A(net439),
    .B(_02913_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02916_));
 sky130_fd_sc_hd__nand2_1 _06003_ (.A(net542),
    .B(net452),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02917_));
 sky130_fd_sc_hd__nor2_1 _06004_ (.A(_02916_),
    .B(_02917_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02918_));
 sky130_fd_sc_hd__a21oi_1 _06005_ (.A1(\top.translation.write_fin ),
    .A2(\top.TRN_sram_complete ),
    .B1(\top.translation.totalEn ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02919_));
 sky130_fd_sc_hd__or4b_1 _06006_ (.A(net441),
    .B(net513),
    .C(_02919_),
    .D_N(_02807_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02920_));
 sky130_fd_sc_hd__a21o_1 _06007_ (.A1(\top.translation.totalEn ),
    .A2(_02814_),
    .B1(_02920_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02921_));
 sky130_fd_sc_hd__inv_2 _06008_ (.A(_02921_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02922_));
 sky130_fd_sc_hd__o21a_1 _06009_ (.A1(_02917_),
    .A2(_02921_),
    .B1(\top.TRN_sram_complete ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02923_));
 sky130_fd_sc_hd__or2_1 _06010_ (.A(net304),
    .B(_02923_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02182_));
 sky130_fd_sc_hd__and3_2 _06011_ (.A(net481),
    .B(\top.controller.state_reg[4] ),
    .C(_02878_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02924_));
 sky130_fd_sc_hd__and3_1 _06012_ (.A(\top.sram_interface.init_counter[1] ),
    .B(\top.sram_interface.init_counter[0] ),
    .C(_02924_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02925_));
 sky130_fd_sc_hd__and3_1 _06013_ (.A(\top.sram_interface.init_counter[2] ),
    .B(\top.sram_interface.init_counter[1] ),
    .C(\top.sram_interface.init_counter[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02926_));
 sky130_fd_sc_hd__and2_1 _06014_ (.A(\top.sram_interface.init_counter[3] ),
    .B(_02926_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02927_));
 sky130_fd_sc_hd__and2_1 _06015_ (.A(_02924_),
    .B(_02927_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02928_));
 sky130_fd_sc_hd__and3_1 _06016_ (.A(\top.sram_interface.init_counter[5] ),
    .B(\top.sram_interface.init_counter[4] ),
    .C(_02928_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02929_));
 sky130_fd_sc_hd__and2_1 _06017_ (.A(\top.sram_interface.init_counter[6] ),
    .B(_02929_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02930_));
 sky130_fd_sc_hd__and3_1 _06018_ (.A(\top.sram_interface.init_counter[8] ),
    .B(\top.sram_interface.init_counter[7] ),
    .C(_02930_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02931_));
 sky130_fd_sc_hd__a31o_1 _06019_ (.A1(\top.sram_interface.init_counter[10] ),
    .A2(\top.sram_interface.init_counter[9] ),
    .A3(_02931_),
    .B1(net1101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02169_));
 sky130_fd_sc_hd__nand2_1 _06020_ (.A(\top.sram_interface.init_counter[9] ),
    .B(_02931_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02932_));
 sky130_fd_sc_hd__xnor2_1 _06021_ (.A(net1518),
    .B(_02932_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02168_));
 sky130_fd_sc_hd__or2_1 _06022_ (.A(\top.sram_interface.init_counter[9] ),
    .B(_02931_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02933_));
 sky130_fd_sc_hd__and2_1 _06023_ (.A(_02932_),
    .B(_02933_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02167_));
 sky130_fd_sc_hd__a21oi_1 _06024_ (.A1(\top.sram_interface.init_counter[7] ),
    .A2(_02930_),
    .B1(\top.sram_interface.init_counter[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02934_));
 sky130_fd_sc_hd__nor2_1 _06025_ (.A(_02931_),
    .B(_02934_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02166_));
 sky130_fd_sc_hd__xor2_1 _06026_ (.A(net1757),
    .B(_02930_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02165_));
 sky130_fd_sc_hd__nor2_1 _06027_ (.A(net1748),
    .B(_02929_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02935_));
 sky130_fd_sc_hd__nor2_1 _06028_ (.A(_02930_),
    .B(_02935_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02164_));
 sky130_fd_sc_hd__a21oi_1 _06029_ (.A1(\top.sram_interface.init_counter[4] ),
    .A2(_02928_),
    .B1(\top.sram_interface.init_counter[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02936_));
 sky130_fd_sc_hd__nor2_1 _06030_ (.A(_02929_),
    .B(_02936_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02163_));
 sky130_fd_sc_hd__xor2_1 _06031_ (.A(net1626),
    .B(_02928_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02162_));
 sky130_fd_sc_hd__a21oi_1 _06032_ (.A1(_02924_),
    .A2(_02926_),
    .B1(net1702),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02937_));
 sky130_fd_sc_hd__nor2_1 _06033_ (.A(_02928_),
    .B(_02937_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02161_));
 sky130_fd_sc_hd__nor2_1 _06034_ (.A(net1614),
    .B(_02925_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02938_));
 sky130_fd_sc_hd__a21oi_1 _06035_ (.A1(_02924_),
    .A2(_02926_),
    .B1(_02938_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02160_));
 sky130_fd_sc_hd__a21oi_1 _06036_ (.A1(\top.sram_interface.init_counter[0] ),
    .A2(_02924_),
    .B1(\top.sram_interface.init_counter[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02939_));
 sky130_fd_sc_hd__nor2_1 _06037_ (.A(_02925_),
    .B(_02939_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02159_));
 sky130_fd_sc_hd__xor2_1 _06038_ (.A(\top.sram_interface.init_counter[0] ),
    .B(_02924_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02158_));
 sky130_fd_sc_hd__or4_1 _06039_ (.A(\top.sram_interface.init_counter[5] ),
    .B(\top.sram_interface.init_counter[4] ),
    .C(\top.sram_interface.init_counter[3] ),
    .D(\top.sram_interface.init_counter[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02940_));
 sky130_fd_sc_hd__or4_1 _06040_ (.A(\top.sram_interface.init_counter[9] ),
    .B(\top.sram_interface.init_counter[8] ),
    .C(\top.sram_interface.init_counter[7] ),
    .D(\top.sram_interface.init_counter[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02941_));
 sky130_fd_sc_hd__or4bb_1 _06041_ (.A(net444),
    .B(\top.sram_interface.init_counter[10] ),
    .C_N(\top.WB.prev_BUSY_O ),
    .D_N(\top.sram_interface.init_counter[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02942_));
 sky130_fd_sc_hd__or4_1 _06042_ (.A(\top.sram_interface.init_counter[1] ),
    .B(\top.sram_interface.init_counter[0] ),
    .C(_02610_),
    .D(_02942_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02943_));
 sky130_fd_sc_hd__or4_1 _06043_ (.A(_02876_),
    .B(_02940_),
    .C(_02941_),
    .D(_02943_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02944_));
 sky130_fd_sc_hd__nand2_1 _06044_ (.A(_02447_),
    .B(_02944_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02157_));
 sky130_fd_sc_hd__a22o_1 _06045_ (.A1(_02449_),
    .A2(\top.cb_syn.zeroes[4] ),
    .B1(\top.cb_syn.zeroes[3] ),
    .B2(_02450_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02945_));
 sky130_fd_sc_hd__o211a_1 _06046_ (.A1(_02452_),
    .A2(\top.cb_syn.zeroes[1] ),
    .B1(\top.cb_syn.zeroes[0] ),
    .C1(_02453_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02946_));
 sky130_fd_sc_hd__a221o_1 _06047_ (.A1(_02451_),
    .A2(\top.cb_syn.zeroes[2] ),
    .B1(\top.cb_syn.zeroes[1] ),
    .B2(_02452_),
    .C1(_02946_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02947_));
 sky130_fd_sc_hd__o22a_1 _06048_ (.A1(_02450_),
    .A2(\top.cb_syn.zeroes[3] ),
    .B1(\top.cb_syn.zeroes[2] ),
    .B2(_02451_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02948_));
 sky130_fd_sc_hd__a21o_1 _06049_ (.A1(_02947_),
    .A2(_02948_),
    .B1(_02945_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02949_));
 sky130_fd_sc_hd__o221a_1 _06050_ (.A1(_02448_),
    .A2(\top.cb_syn.zeroes[5] ),
    .B1(\top.cb_syn.zeroes[4] ),
    .B2(_02449_),
    .C1(_02949_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02950_));
 sky130_fd_sc_hd__nor2_1 _06051_ (.A(\top.cb_syn.count[5] ),
    .B(_02528_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02951_));
 sky130_fd_sc_hd__a2bb2o_1 _06052_ (.A1_N(_02950_),
    .A2_N(_02951_),
    .B1(\top.cb_syn.count[6] ),
    .B2(_02527_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02952_));
 sky130_fd_sc_hd__o221a_1 _06053_ (.A1(\top.cb_syn.count[7] ),
    .A2(_02526_),
    .B1(_02527_),
    .B2(\top.cb_syn.count[6] ),
    .C1(_02952_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02953_));
 sky130_fd_sc_hd__a22o_1 _06054_ (.A1(_02528_),
    .A2(\top.cb_syn.zero_count[5] ),
    .B1(\top.cb_syn.zero_count[4] ),
    .B2(_02529_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02954_));
 sky130_fd_sc_hd__nand2_1 _06055_ (.A(_02527_),
    .B(\top.cb_syn.zero_count[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02955_));
 sky130_fd_sc_hd__a22o_1 _06056_ (.A1(_02533_),
    .A2(\top.cb_syn.zero_count[0] ),
    .B1(\top.cb_syn.zero_count[1] ),
    .B2(_02532_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02956_));
 sky130_fd_sc_hd__a2bb2o_1 _06057_ (.A1_N(_02527_),
    .A2_N(\top.cb_syn.zero_count[6] ),
    .B1(_02559_),
    .B2(\top.cb_syn.zeroes[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02957_));
 sky130_fd_sc_hd__o22a_1 _06058_ (.A1(_02530_),
    .A2(\top.cb_syn.zero_count[3] ),
    .B1(\top.cb_syn.zero_count[2] ),
    .B2(_02531_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02958_));
 sky130_fd_sc_hd__nor2_1 _06059_ (.A(\top.cb_syn.zeroes[3] ),
    .B(_02557_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02959_));
 sky130_fd_sc_hd__nor2_1 _06060_ (.A(\top.cb_syn.zeroes[2] ),
    .B(_02558_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02960_));
 sky130_fd_sc_hd__or3b_1 _06061_ (.A(_02959_),
    .B(_02960_),
    .C_N(_02958_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02961_));
 sky130_fd_sc_hd__nor2_1 _06062_ (.A(_02526_),
    .B(\top.cb_syn.zero_count[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02962_));
 sky130_fd_sc_hd__and2_1 _06063_ (.A(_02526_),
    .B(\top.cb_syn.zero_count[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02963_));
 sky130_fd_sc_hd__or2_1 _06064_ (.A(_02532_),
    .B(\top.cb_syn.zero_count[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02964_));
 sky130_fd_sc_hd__o211a_1 _06065_ (.A1(_02529_),
    .A2(\top.cb_syn.zero_count[4] ),
    .B1(_02955_),
    .C1(_02964_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02965_));
 sky130_fd_sc_hd__a211o_1 _06066_ (.A1(\top.cb_syn.zeroes[0] ),
    .A2(_02556_),
    .B1(_02956_),
    .C1(_02962_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02966_));
 sky130_fd_sc_hd__or4_1 _06067_ (.A(_02954_),
    .B(_02957_),
    .C(_02961_),
    .D(_02966_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02967_));
 sky130_fd_sc_hd__nor3b_1 _06068_ (.A(_02967_),
    .B(_02963_),
    .C_N(_02965_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02968_));
 sky130_fd_sc_hd__a211oi_2 _06069_ (.A1(\top.cb_syn.count[7] ),
    .A2(_02526_),
    .B1(_02953_),
    .C1(_02968_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02969_));
 sky130_fd_sc_hd__nand2b_1 _06070_ (.A_N(\top.cb_syn.cb_length[6] ),
    .B(\top.cb_syn.i[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02970_));
 sky130_fd_sc_hd__nand2b_1 _06071_ (.A_N(\top.cb_syn.i[6] ),
    .B(\top.cb_syn.cb_length[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02971_));
 sky130_fd_sc_hd__nand2_1 _06072_ (.A(_02970_),
    .B(_02971_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02972_));
 sky130_fd_sc_hd__and2b_1 _06073_ (.A_N(\top.cb_syn.cb_length[2] ),
    .B(\top.cb_syn.i[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02973_));
 sky130_fd_sc_hd__and2b_1 _06074_ (.A_N(\top.cb_syn.i[2] ),
    .B(\top.cb_syn.cb_length[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02974_));
 sky130_fd_sc_hd__nor2_2 _06075_ (.A(_02973_),
    .B(_02974_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02975_));
 sky130_fd_sc_hd__inv_2 _06076_ (.A(_02975_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02976_));
 sky130_fd_sc_hd__nand2_1 _06077_ (.A(_02534_),
    .B(\top.cb_syn.i[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02977_));
 sky130_fd_sc_hd__or2_1 _06078_ (.A(_02534_),
    .B(\top.cb_syn.i[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02978_));
 sky130_fd_sc_hd__nand2_2 _06079_ (.A(_02977_),
    .B(_02978_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02979_));
 sky130_fd_sc_hd__nand2b_1 _06080_ (.A_N(\top.cb_syn.cb_length[0] ),
    .B(\top.cb_syn.i[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02980_));
 sky130_fd_sc_hd__xnor2_1 _06081_ (.A(\top.cb_syn.cb_length[0] ),
    .B(\top.cb_syn.i[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02981_));
 sky130_fd_sc_hd__and2b_1 _06082_ (.A_N(\top.cb_syn.i[1] ),
    .B(\top.cb_syn.cb_length[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02982_));
 sky130_fd_sc_hd__and2b_1 _06083_ (.A_N(\top.cb_syn.cb_length[1] ),
    .B(\top.cb_syn.i[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02983_));
 sky130_fd_sc_hd__nor2_1 _06084_ (.A(_02982_),
    .B(_02983_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02984_));
 sky130_fd_sc_hd__and2b_1 _06085_ (.A_N(\top.cb_syn.cb_length[5] ),
    .B(\top.cb_syn.i[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02985_));
 sky130_fd_sc_hd__and2b_1 _06086_ (.A_N(\top.cb_syn.i[5] ),
    .B(\top.cb_syn.cb_length[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02986_));
 sky130_fd_sc_hd__or2_1 _06087_ (.A(_02985_),
    .B(_02986_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02987_));
 sky130_fd_sc_hd__inv_2 _06088_ (.A(_02987_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02988_));
 sky130_fd_sc_hd__and2_1 _06089_ (.A(_02535_),
    .B(\top.cb_syn.i[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02989_));
 sky130_fd_sc_hd__nor2_1 _06090_ (.A(_02535_),
    .B(\top.cb_syn.i[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02990_));
 sky130_fd_sc_hd__or2_2 _06091_ (.A(_02989_),
    .B(_02990_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02991_));
 sky130_fd_sc_hd__nor4_1 _06092_ (.A(_02972_),
    .B(_02976_),
    .C(_02987_),
    .D(_02991_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02992_));
 sky130_fd_sc_hd__and4b_1 _06093_ (.A_N(_02979_),
    .B(net394),
    .C(_02984_),
    .D(_02992_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02993_));
 sky130_fd_sc_hd__nor2_1 _06094_ (.A(_02969_),
    .B(_02993_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02994_));
 sky130_fd_sc_hd__and2_1 _06095_ (.A(net550),
    .B(_02994_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02995_));
 sky130_fd_sc_hd__or3_4 _06096_ (.A(_02554_),
    .B(net423),
    .C(_02995_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02996_));
 sky130_fd_sc_hd__and3_2 _06097_ (.A(net523),
    .B(net463),
    .C(_02969_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02997_));
 sky130_fd_sc_hd__nand2_1 _06098_ (.A(\top.cb_syn.count[1] ),
    .B(\top.cb_syn.count[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02998_));
 sky130_fd_sc_hd__or2_1 _06099_ (.A(_02451_),
    .B(_02998_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02999_));
 sky130_fd_sc_hd__nor2_1 _06100_ (.A(_02450_),
    .B(_02999_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03000_));
 sky130_fd_sc_hd__inv_2 _06101_ (.A(_03000_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03001_));
 sky130_fd_sc_hd__nand2_1 _06102_ (.A(\top.cb_syn.count[4] ),
    .B(_03000_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03002_));
 sky130_fd_sc_hd__nor2_1 _06103_ (.A(_02448_),
    .B(_03002_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03003_));
 sky130_fd_sc_hd__inv_2 _06104_ (.A(_03003_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03004_));
 sky130_fd_sc_hd__nand2_1 _06105_ (.A(\top.cb_syn.count[6] ),
    .B(_03003_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03005_));
 sky130_fd_sc_hd__xnor2_1 _06106_ (.A(\top.cb_syn.count[7] ),
    .B(_03005_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03006_));
 sky130_fd_sc_hd__a22o_1 _06107_ (.A1(\top.cb_syn.count[7] ),
    .A2(_02996_),
    .B1(_02997_),
    .B2(_03006_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02156_));
 sky130_fd_sc_hd__or2_1 _06108_ (.A(\top.cb_syn.count[6] ),
    .B(_03003_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03007_));
 sky130_fd_sc_hd__a32o_1 _06109_ (.A1(_02997_),
    .A2(_03005_),
    .A3(_03007_),
    .B1(_02996_),
    .B2(net1641),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02155_));
 sky130_fd_sc_hd__nand2_1 _06110_ (.A(_02448_),
    .B(_03002_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03008_));
 sky130_fd_sc_hd__a32o_1 _06111_ (.A1(_02997_),
    .A2(_03004_),
    .A3(_03008_),
    .B1(_02996_),
    .B2(net1595),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02154_));
 sky130_fd_sc_hd__or2_1 _06112_ (.A(\top.cb_syn.count[4] ),
    .B(_03000_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03009_));
 sky130_fd_sc_hd__a32o_1 _06113_ (.A1(_02997_),
    .A2(_03002_),
    .A3(_03009_),
    .B1(_02996_),
    .B2(net1662),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02153_));
 sky130_fd_sc_hd__nand2_1 _06114_ (.A(_02450_),
    .B(_02999_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03010_));
 sky130_fd_sc_hd__a32o_1 _06115_ (.A1(_02997_),
    .A2(_03001_),
    .A3(_03010_),
    .B1(_02996_),
    .B2(net1438),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02152_));
 sky130_fd_sc_hd__nand2_1 _06116_ (.A(_02451_),
    .B(_02998_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03011_));
 sky130_fd_sc_hd__a32o_1 _06117_ (.A1(_02997_),
    .A2(_02999_),
    .A3(_03011_),
    .B1(_02996_),
    .B2(net1463),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02151_));
 sky130_fd_sc_hd__or2_1 _06118_ (.A(\top.cb_syn.count[1] ),
    .B(\top.cb_syn.count[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03012_));
 sky130_fd_sc_hd__a32o_1 _06119_ (.A1(_02997_),
    .A2(_02998_),
    .A3(_03012_),
    .B1(_02996_),
    .B2(net1673),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02150_));
 sky130_fd_sc_hd__mux2_1 _06120_ (.A0(_02996_),
    .A1(_02997_),
    .S(_02453_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02149_));
 sky130_fd_sc_hd__a31o_1 _06121_ (.A1(net453),
    .A2(\top.histogram.eof_n ),
    .A3(_02561_),
    .B1(net1034),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02148_));
 sky130_fd_sc_hd__a21o_1 _06122_ (.A1(net1434),
    .A2(_02619_),
    .B1(net207),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02147_));
 sky130_fd_sc_hd__and2_1 _06123_ (.A(net1053),
    .B(net166),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02146_));
 sky130_fd_sc_hd__a21o_1 _06124_ (.A1(net1018),
    .A2(_02619_),
    .B1(net207),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02145_));
 sky130_fd_sc_hd__or2_2 _06125_ (.A(net461),
    .B(\top.controller.state_reg[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03013_));
 sky130_fd_sc_hd__o21ai_1 _06126_ (.A1(net542),
    .A2(net526),
    .B1(net406),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03014_));
 sky130_fd_sc_hd__or4_1 _06127_ (.A(net444),
    .B(net453),
    .C(net447),
    .D(_03014_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03015_));
 sky130_fd_sc_hd__or4_1 _06128_ (.A(net533),
    .B(net527),
    .C(_03013_),
    .D(_03015_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03016_));
 sky130_fd_sc_hd__a22o_1 _06129_ (.A1(net1226),
    .A2(net164),
    .B1(_03016_),
    .B2(net207),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02144_));
 sky130_fd_sc_hd__and4_2 _06130_ (.A(net458),
    .B(net361),
    .C(net208),
    .D(net407),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03017_));
 sky130_fd_sc_hd__a21o_1 _06131_ (.A1(net1466),
    .A2(net164),
    .B1(net157),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02143_));
 sky130_fd_sc_hd__a21o_1 _06132_ (.A1(net1036),
    .A2(net166),
    .B1(net157),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02142_));
 sky130_fd_sc_hd__a21o_1 _06133_ (.A1(net1033),
    .A2(net166),
    .B1(net157),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02141_));
 sky130_fd_sc_hd__a21o_1 _06134_ (.A1(net1012),
    .A2(net166),
    .B1(net157),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02140_));
 sky130_fd_sc_hd__a21o_1 _06135_ (.A1(net1042),
    .A2(net166),
    .B1(net157),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02139_));
 sky130_fd_sc_hd__a21o_1 _06136_ (.A1(net1031),
    .A2(net166),
    .B1(net157),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02138_));
 sky130_fd_sc_hd__a21o_1 _06137_ (.A1(net1587),
    .A2(net164),
    .B1(net157),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02137_));
 sky130_fd_sc_hd__a21o_1 _06138_ (.A1(net1043),
    .A2(net166),
    .B1(net157),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02136_));
 sky130_fd_sc_hd__a21o_1 _06139_ (.A1(net1032),
    .A2(net166),
    .B1(_03017_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02135_));
 sky130_fd_sc_hd__a21o_1 _06140_ (.A1(net1093),
    .A2(net166),
    .B1(_03017_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02134_));
 sky130_fd_sc_hd__and2_1 _06141_ (.A(net481),
    .B(_02877_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03018_));
 sky130_fd_sc_hd__nand2_2 _06142_ (.A(net481),
    .B(_02877_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03019_));
 sky130_fd_sc_hd__nor2_1 _06143_ (.A(\top.sram_interface.init_counter[3] ),
    .B(_02926_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03020_));
 sky130_fd_sc_hd__o21a_1 _06144_ (.A1(\top.sram_interface.init_counter[3] ),
    .A2(_02926_),
    .B1(\top.sram_interface.init_counter[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03021_));
 sky130_fd_sc_hd__and2_1 _06145_ (.A(\top.sram_interface.init_counter[5] ),
    .B(_03021_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03022_));
 sky130_fd_sc_hd__and3_1 _06146_ (.A(\top.sram_interface.init_counter[6] ),
    .B(\top.sram_interface.init_counter[5] ),
    .C(_03021_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03023_));
 sky130_fd_sc_hd__and3_1 _06147_ (.A(\top.sram_interface.init_counter[8] ),
    .B(\top.sram_interface.init_counter[7] ),
    .C(_03023_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03024_));
 sky130_fd_sc_hd__and2_1 _06148_ (.A(\top.sram_interface.init_counter[9] ),
    .B(_03024_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03025_));
 sky130_fd_sc_hd__o21ai_1 _06149_ (.A1(\top.sram_interface.init_counter[10] ),
    .A2(_03025_),
    .B1(_03018_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03026_));
 sky130_fd_sc_hd__nor3b_1 _06150_ (.A(_02417_),
    .B(_03026_),
    .C_N(net207),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03027_));
 sky130_fd_sc_hd__a211o_1 _06151_ (.A1(net1048),
    .A2(net164),
    .B1(net157),
    .C1(_03027_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02133_));
 sky130_fd_sc_hd__a21o_1 _06152_ (.A1(\top.sram_interface.init_counter[10] ),
    .A2(_03025_),
    .B1(_03026_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03028_));
 sky130_fd_sc_hd__a31o_1 _06153_ (.A1(net458),
    .A2(net533),
    .A3(net407),
    .B1(_02592_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03029_));
 sky130_fd_sc_hd__a211o_1 _06154_ (.A1(net454),
    .A2(_03028_),
    .B1(_03029_),
    .C1(_02608_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03030_));
 sky130_fd_sc_hd__a221o_1 _06155_ (.A1(net1525),
    .A2(net164),
    .B1(_03030_),
    .B2(net207),
    .C1(net157),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02132_));
 sky130_fd_sc_hd__nor2_1 _06156_ (.A(\top.sram_interface.init_counter[9] ),
    .B(_03024_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03031_));
 sky130_fd_sc_hd__o21a_1 _06157_ (.A1(_03025_),
    .A2(_03031_),
    .B1(_02877_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03032_));
 sky130_fd_sc_hd__nor2_1 _06158_ (.A(_02610_),
    .B(_03032_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03033_));
 sky130_fd_sc_hd__nand2_1 _06159_ (.A(\top.cb_syn.char_index[2] ),
    .B(\top.cb_syn.char_index[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03034_));
 sky130_fd_sc_hd__and4_1 _06160_ (.A(\top.cb_syn.char_index[4] ),
    .B(\top.cb_syn.char_index[3] ),
    .C(\top.cb_syn.char_index[2] ),
    .D(\top.cb_syn.char_index[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03035_));
 sky130_fd_sc_hd__nand2_1 _06161_ (.A(\top.cb_syn.char_index[5] ),
    .B(_03035_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03036_));
 sky130_fd_sc_hd__nand2_1 _06162_ (.A(\top.findLeastValue.histo_index[8] ),
    .B(\top.findLeastValue.histo_index[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03037_));
 sky130_fd_sc_hd__and3_1 _06163_ (.A(net459),
    .B(net534),
    .C(_02787_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03038_));
 sky130_fd_sc_hd__a21oi_1 _06164_ (.A1(net459),
    .A2(net361),
    .B1(_03038_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03039_));
 sky130_fd_sc_hd__a21oi_1 _06165_ (.A1(_02787_),
    .A2(_03037_),
    .B1(_03039_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03040_));
 sky130_fd_sc_hd__a41o_1 _06166_ (.A1(\top.cb_syn.char_index[6] ),
    .A2(\top.cb_syn.char_index[5] ),
    .A3(_02607_),
    .A4(_03035_),
    .B1(_03040_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03041_));
 sky130_fd_sc_hd__or2_1 _06167_ (.A(\top.cb_syn.char_index[1] ),
    .B(\top.cb_syn.char_index[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03042_));
 sky130_fd_sc_hd__nand2_1 _06168_ (.A(\top.cb_syn.char_index[2] ),
    .B(_03042_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03043_));
 sky130_fd_sc_hd__and3_1 _06169_ (.A(\top.cb_syn.char_index[3] ),
    .B(\top.cb_syn.char_index[2] ),
    .C(_03042_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03044_));
 sky130_fd_sc_hd__inv_2 _06170_ (.A(_03044_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03045_));
 sky130_fd_sc_hd__and2_1 _06171_ (.A(\top.cb_syn.char_index[4] ),
    .B(_03044_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03046_));
 sky130_fd_sc_hd__and3_1 _06172_ (.A(\top.cb_syn.char_index[5] ),
    .B(\top.cb_syn.char_index[4] ),
    .C(_03044_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03047_));
 sky130_fd_sc_hd__or3b_1 _06173_ (.A(_02536_),
    .B(_02605_),
    .C_N(_03047_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03048_));
 sky130_fd_sc_hd__nand2_1 _06174_ (.A(net445),
    .B(\top.TRN_char_index[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03049_));
 sky130_fd_sc_hd__and3_1 _06175_ (.A(\top.TRN_char_index[3] ),
    .B(net445),
    .C(\top.TRN_char_index[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03050_));
 sky130_fd_sc_hd__and3_1 _06176_ (.A(\top.TRN_char_index[5] ),
    .B(\top.TRN_char_index[4] ),
    .C(_03050_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03051_));
 sky130_fd_sc_hd__nand2_1 _06177_ (.A(\top.TRN_char_index[6] ),
    .B(_03051_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03052_));
 sky130_fd_sc_hd__or2_1 _06178_ (.A(\top.TRN_char_index[1] ),
    .B(\top.TRN_char_index[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03053_));
 sky130_fd_sc_hd__nand2_1 _06179_ (.A(net445),
    .B(_03053_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03054_));
 sky130_fd_sc_hd__and3_1 _06180_ (.A(\top.TRN_char_index[3] ),
    .B(net445),
    .C(_03053_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03055_));
 sky130_fd_sc_hd__and2_1 _06181_ (.A(\top.TRN_char_index[4] ),
    .B(_03055_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03056_));
 sky130_fd_sc_hd__and3_1 _06182_ (.A(\top.TRN_char_index[5] ),
    .B(\top.TRN_char_index[4] ),
    .C(_03055_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03057_));
 sky130_fd_sc_hd__and2_1 _06183_ (.A(net545),
    .B(_03057_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03058_));
 sky130_fd_sc_hd__o211a_1 _06184_ (.A1(_03051_),
    .A2(_03058_),
    .B1(\top.TRN_char_index[6] ),
    .C1(_02592_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03059_));
 sky130_fd_sc_hd__or4b_1 _06185_ (.A(_03033_),
    .B(_03059_),
    .C(_03041_),
    .D_N(_03048_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03060_));
 sky130_fd_sc_hd__a22o_1 _06186_ (.A1(net1548),
    .A2(net164),
    .B1(_03060_),
    .B2(net207),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02131_));
 sky130_fd_sc_hd__a21oi_1 _06187_ (.A1(\top.sram_interface.init_counter[7] ),
    .A2(_03023_),
    .B1(\top.sram_interface.init_counter[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03061_));
 sky130_fd_sc_hd__o21a_1 _06188_ (.A1(_03024_),
    .A2(_03061_),
    .B1(_02877_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03062_));
 sky130_fd_sc_hd__a21oi_1 _06189_ (.A1(\top.cb_syn.char_index[6] ),
    .A2(_03047_),
    .B1(_02605_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03063_));
 sky130_fd_sc_hd__o21a_1 _06190_ (.A1(\top.cb_syn.char_index[6] ),
    .A2(_03047_),
    .B1(_03063_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03064_));
 sky130_fd_sc_hd__a21oi_1 _06191_ (.A1(\top.TRN_char_index[6] ),
    .A2(_03057_),
    .B1(_02585_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03065_));
 sky130_fd_sc_hd__o21a_1 _06192_ (.A1(\top.TRN_char_index[6] ),
    .A2(_03057_),
    .B1(_03065_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03066_));
 sky130_fd_sc_hd__or2_1 _06193_ (.A(\top.TRN_char_index[6] ),
    .B(_03051_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03067_));
 sky130_fd_sc_hd__xnor2_1 _06194_ (.A(\top.cb_syn.char_index[6] ),
    .B(_03036_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03068_));
 sky130_fd_sc_hd__a32o_1 _06195_ (.A1(_02590_),
    .A2(_03052_),
    .A3(_03067_),
    .B1(_03068_),
    .B2(_02607_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03069_));
 sky130_fd_sc_hd__and3_1 _06196_ (.A(\top.cw1[2] ),
    .B(\top.cw1[1] ),
    .C(\top.cw1[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03070_));
 sky130_fd_sc_hd__or2_1 _06197_ (.A(\top.cw1[3] ),
    .B(_03070_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03071_));
 sky130_fd_sc_hd__and3_1 _06198_ (.A(\top.cw1[5] ),
    .B(\top.cw1[4] ),
    .C(_03071_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03072_));
 sky130_fd_sc_hd__and2_1 _06199_ (.A(\top.cw1[6] ),
    .B(_03072_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03073_));
 sky130_fd_sc_hd__a21o_1 _06200_ (.A1(\top.cw1[7] ),
    .A2(_03073_),
    .B1(_02602_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03074_));
 sky130_fd_sc_hd__a41o_1 _06201_ (.A1(\top.findLeastValue.histo_index[8] ),
    .A2(_02501_),
    .A3(net534),
    .A4(_02575_),
    .B1(_02603_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03075_));
 sky130_fd_sc_hd__nand2_1 _06202_ (.A(\top.cw2[1] ),
    .B(\top.cw2[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03076_));
 sky130_fd_sc_hd__nor2_1 _06203_ (.A(_02510_),
    .B(_03076_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03077_));
 sky130_fd_sc_hd__inv_2 _06204_ (.A(_03077_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03078_));
 sky130_fd_sc_hd__o21ai_1 _06205_ (.A1(\top.cw2[3] ),
    .A2(_03077_),
    .B1(\top.cw2[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03079_));
 sky130_fd_sc_hd__nor2_1 _06206_ (.A(_02507_),
    .B(_03079_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03080_));
 sky130_fd_sc_hd__and2_1 _06207_ (.A(\top.cw2[6] ),
    .B(_03080_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03081_));
 sky130_fd_sc_hd__a22o_1 _06208_ (.A1(_02501_),
    .A2(net361),
    .B1(_03074_),
    .B2(_03075_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03082_));
 sky130_fd_sc_hd__a31o_1 _06209_ (.A1(\top.cw2[7] ),
    .A2(_02600_),
    .A3(_03081_),
    .B1(_03082_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03083_));
 sky130_fd_sc_hd__a2bb2o_1 _06210_ (.A1_N(_02610_),
    .A2_N(_03062_),
    .B1(_03083_),
    .B2(net458),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03084_));
 sky130_fd_sc_hd__or4_1 _06211_ (.A(_03064_),
    .B(_03066_),
    .C(_03069_),
    .D(_03084_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03085_));
 sky130_fd_sc_hd__a22o_1 _06212_ (.A1(net1691),
    .A2(net164),
    .B1(_03085_),
    .B2(net208),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02130_));
 sky130_fd_sc_hd__xor2_1 _06213_ (.A(\top.cw1[7] ),
    .B(_03073_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03086_));
 sky130_fd_sc_hd__nand2_1 _06214_ (.A(net487),
    .B(\top.findLeastValue.histo_index[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03087_));
 sky130_fd_sc_hd__and3_1 _06215_ (.A(\top.findLeastValue.histo_index[2] ),
    .B(net487),
    .C(\top.findLeastValue.histo_index[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03088_));
 sky130_fd_sc_hd__or2_2 _06216_ (.A(net486),
    .B(_03088_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03089_));
 sky130_fd_sc_hd__a21oi_1 _06217_ (.A1(net484),
    .A2(_03089_),
    .B1(_02787_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03090_));
 sky130_fd_sc_hd__a31o_1 _06218_ (.A1(net483),
    .A2(net484),
    .A3(_03089_),
    .B1(_02787_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03091_));
 sky130_fd_sc_hd__and3_1 _06219_ (.A(net482),
    .B(net534),
    .C(_03091_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03092_));
 sky130_fd_sc_hd__o22a_1 _06220_ (.A1(_02602_),
    .A2(_03086_),
    .B1(_03092_),
    .B2(_02603_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03093_));
 sky130_fd_sc_hd__xnor2_1 _06221_ (.A(_02505_),
    .B(_03081_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03094_));
 sky130_fd_sc_hd__a221o_1 _06222_ (.A1(net482),
    .A2(net361),
    .B1(_02600_),
    .B2(_03094_),
    .C1(_03093_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03095_));
 sky130_fd_sc_hd__xor2_1 _06223_ (.A(\top.sram_interface.init_counter[7] ),
    .B(_03023_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03096_));
 sky130_fd_sc_hd__nand2_1 _06224_ (.A(\top.hist_addr[1] ),
    .B(\top.hist_addr[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03097_));
 sky130_fd_sc_hd__a31o_1 _06225_ (.A1(\top.hist_addr[2] ),
    .A2(\top.hist_addr[1] ),
    .A3(\top.hist_addr[0] ),
    .B1(\top.hist_addr[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03098_));
 sky130_fd_sc_hd__and3_1 _06226_ (.A(\top.hist_addr[5] ),
    .B(\top.hist_addr[4] ),
    .C(_03098_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03099_));
 sky130_fd_sc_hd__a21o_1 _06227_ (.A1(\top.hist_addr[6] ),
    .A2(_03099_),
    .B1(net481),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03100_));
 sky130_fd_sc_hd__o211a_1 _06228_ (.A1(_03019_),
    .A2(_03096_),
    .B1(_03100_),
    .C1(net454),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03101_));
 sky130_fd_sc_hd__a31o_2 _06229_ (.A1(_02418_),
    .A2(_02524_),
    .A3(net533),
    .B1(\top.sram_interface.word_cnt[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03102_));
 sky130_fd_sc_hd__o21a_1 _06230_ (.A1(\top.hTree.write_HT_fin ),
    .A2(\top.WorR ),
    .B1(net533),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03103_));
 sky130_fd_sc_hd__or3_4 _06231_ (.A(net526),
    .B(\top.sram_interface.word_cnt[13] ),
    .C(_03103_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03104_));
 sky130_fd_sc_hd__a22o_1 _06232_ (.A1(\top.cb_syn.max_index[7] ),
    .A2(_03102_),
    .B1(_03104_),
    .B2(\top.hTree.nullSumIndex[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03105_));
 sky130_fd_sc_hd__nor2_1 _06233_ (.A(_02585_),
    .B(_03057_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03106_));
 sky130_fd_sc_hd__o21a_1 _06234_ (.A1(\top.TRN_char_index[5] ),
    .A2(_03056_),
    .B1(_03106_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03107_));
 sky130_fd_sc_hd__a21oi_1 _06235_ (.A1(\top.TRN_char_index[4] ),
    .A2(_03050_),
    .B1(\top.TRN_char_index[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03108_));
 sky130_fd_sc_hd__nor3_1 _06236_ (.A(_02591_),
    .B(_03051_),
    .C(_03108_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03109_));
 sky130_fd_sc_hd__nor2_1 _06237_ (.A(_02605_),
    .B(_03047_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03110_));
 sky130_fd_sc_hd__o21a_1 _06238_ (.A1(\top.cb_syn.char_index[5] ),
    .A2(_03046_),
    .B1(_03110_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03111_));
 sky130_fd_sc_hd__or2_1 _06239_ (.A(\top.cb_syn.char_index[5] ),
    .B(_03035_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03112_));
 sky130_fd_sc_hd__a22o_1 _06240_ (.A1(\top.cb_syn.curr_index[7] ),
    .A2(_02584_),
    .B1(_03105_),
    .B2(net446),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03113_));
 sky130_fd_sc_hd__a31o_1 _06241_ (.A1(_02607_),
    .A2(_03036_),
    .A3(_03112_),
    .B1(_03107_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03114_));
 sky130_fd_sc_hd__or4_1 _06242_ (.A(_03109_),
    .B(_03111_),
    .C(_03113_),
    .D(_03114_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03115_));
 sky130_fd_sc_hd__a211o_1 _06243_ (.A1(net458),
    .A2(_03095_),
    .B1(_03101_),
    .C1(_03115_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03116_));
 sky130_fd_sc_hd__a22o_1 _06244_ (.A1(net1379),
    .A2(net164),
    .B1(_03116_),
    .B2(net207),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02129_));
 sky130_fd_sc_hd__nor2_1 _06245_ (.A(\top.cw1[6] ),
    .B(_03072_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03117_));
 sky130_fd_sc_hd__or2_1 _06246_ (.A(\top.cw2[6] ),
    .B(_03080_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03118_));
 sky130_fd_sc_hd__and3b_1 _06247_ (.A_N(_03081_),
    .B(_03118_),
    .C(_02600_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03119_));
 sky130_fd_sc_hd__a211o_1 _06248_ (.A1(net482),
    .A2(net406),
    .B1(_03090_),
    .C1(_02503_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03120_));
 sky130_fd_sc_hd__o31a_1 _06249_ (.A1(_02602_),
    .A2(_03073_),
    .A3(_03117_),
    .B1(_03120_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03121_));
 sky130_fd_sc_hd__o21ai_1 _06250_ (.A1(_02502_),
    .A2(_03091_),
    .B1(_03121_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03122_));
 sky130_fd_sc_hd__a22o_1 _06251_ (.A1(net483),
    .A2(net361),
    .B1(_03122_),
    .B2(net534),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03123_));
 sky130_fd_sc_hd__o21a_1 _06252_ (.A1(_03119_),
    .A2(_03123_),
    .B1(net459),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03124_));
 sky130_fd_sc_hd__xor2_1 _06253_ (.A(\top.hist_addr[6] ),
    .B(_03099_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03125_));
 sky130_fd_sc_hd__nor2_1 _06254_ (.A(\top.sram_interface.init_counter[6] ),
    .B(_03022_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03126_));
 sky130_fd_sc_hd__nor2_1 _06255_ (.A(_03023_),
    .B(_03126_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03127_));
 sky130_fd_sc_hd__o221a_1 _06256_ (.A1(net481),
    .A2(_03125_),
    .B1(_03127_),
    .B2(_03019_),
    .C1(net454),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03128_));
 sky130_fd_sc_hd__a31o_1 _06257_ (.A1(\top.cb_syn.char_index[3] ),
    .A2(\top.cb_syn.char_index[2] ),
    .A3(\top.cb_syn.char_index[1] ),
    .B1(\top.cb_syn.char_index[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03129_));
 sky130_fd_sc_hd__and3b_1 _06258_ (.A_N(_03035_),
    .B(_03129_),
    .C(_02607_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03130_));
 sky130_fd_sc_hd__nor2_1 _06259_ (.A(\top.TRN_char_index[4] ),
    .B(_03055_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03131_));
 sky130_fd_sc_hd__a21oi_1 _06260_ (.A1(\top.TRN_char_index[4] ),
    .A2(_03050_),
    .B1(_02591_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03132_));
 sky130_fd_sc_hd__o21ai_1 _06261_ (.A1(\top.TRN_char_index[4] ),
    .A2(_03050_),
    .B1(_03132_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03133_));
 sky130_fd_sc_hd__a22o_1 _06262_ (.A1(\top.cb_syn.max_index[6] ),
    .A2(_03102_),
    .B1(_03104_),
    .B2(\top.hTree.nullSumIndex[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03134_));
 sky130_fd_sc_hd__nor2_1 _06263_ (.A(\top.cb_syn.char_index[4] ),
    .B(_03044_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03135_));
 sky130_fd_sc_hd__or3_1 _06264_ (.A(_02605_),
    .B(_03046_),
    .C(_03135_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03136_));
 sky130_fd_sc_hd__o311a_1 _06265_ (.A1(_02585_),
    .A2(_03056_),
    .A3(_03131_),
    .B1(_03133_),
    .C1(_03136_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03137_));
 sky130_fd_sc_hd__a221o_1 _06266_ (.A1(\top.cb_syn.curr_index[6] ),
    .A2(_02584_),
    .B1(_03134_),
    .B2(net446),
    .C1(_03130_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03138_));
 sky130_fd_sc_hd__or4b_1 _06267_ (.A(_03124_),
    .B(_03138_),
    .C(_03128_),
    .D_N(_03137_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03139_));
 sky130_fd_sc_hd__a22o_1 _06268_ (.A1(net1233),
    .A2(net164),
    .B1(_03139_),
    .B2(net207),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02128_));
 sky130_fd_sc_hd__a21oi_1 _06269_ (.A1(net484),
    .A2(_03089_),
    .B1(net483),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03140_));
 sky130_fd_sc_hd__a2bb2o_1 _06270_ (.A1_N(_03091_),
    .A2_N(_03140_),
    .B1(net484),
    .B2(_02787_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03141_));
 sky130_fd_sc_hd__a21oi_1 _06271_ (.A1(\top.cw1[4] ),
    .A2(_03071_),
    .B1(\top.cw1[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03142_));
 sky130_fd_sc_hd__o21ai_1 _06272_ (.A1(_03072_),
    .A2(_03142_),
    .B1(_02601_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03143_));
 sky130_fd_sc_hd__o211a_1 _06273_ (.A1(_02601_),
    .A2(_03141_),
    .B1(_03143_),
    .C1(net534),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03144_));
 sky130_fd_sc_hd__nand2_1 _06274_ (.A(_02507_),
    .B(_03079_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03145_));
 sky130_fd_sc_hd__and3b_1 _06275_ (.A_N(_03080_),
    .B(_03145_),
    .C(_02600_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03146_));
 sky130_fd_sc_hd__a211o_1 _06276_ (.A1(net484),
    .A2(net361),
    .B1(_03144_),
    .C1(_03146_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03147_));
 sky130_fd_sc_hd__a21oi_1 _06277_ (.A1(\top.hist_addr[4] ),
    .A2(_03098_),
    .B1(\top.hist_addr[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03148_));
 sky130_fd_sc_hd__o21ai_1 _06278_ (.A1(_03099_),
    .A2(_03148_),
    .B1(_02416_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03149_));
 sky130_fd_sc_hd__nor2_1 _06279_ (.A(\top.sram_interface.init_counter[5] ),
    .B(_03021_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03150_));
 sky130_fd_sc_hd__o21ai_1 _06280_ (.A1(_03022_),
    .A2(_03150_),
    .B1(_03018_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03151_));
 sky130_fd_sc_hd__xnor2_1 _06281_ (.A(\top.cb_syn.char_index[3] ),
    .B(_03034_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03152_));
 sky130_fd_sc_hd__a22o_1 _06282_ (.A1(\top.cb_syn.max_index[5] ),
    .A2(_03102_),
    .B1(_03104_),
    .B2(\top.hTree.nullSumIndex[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03153_));
 sky130_fd_sc_hd__nand2_1 _06283_ (.A(net446),
    .B(_03153_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03154_));
 sky130_fd_sc_hd__a21oi_1 _06284_ (.A1(net445),
    .A2(_03053_),
    .B1(\top.TRN_char_index[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03155_));
 sky130_fd_sc_hd__a21oi_1 _06285_ (.A1(net445),
    .A2(\top.TRN_char_index[1] ),
    .B1(\top.TRN_char_index[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03156_));
 sky130_fd_sc_hd__or3_1 _06286_ (.A(_02591_),
    .B(_03050_),
    .C(_03156_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03157_));
 sky130_fd_sc_hd__o311a_1 _06287_ (.A1(_02585_),
    .A2(_03055_),
    .A3(_03155_),
    .B1(_03157_),
    .C1(_03154_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03158_));
 sky130_fd_sc_hd__a21o_1 _06288_ (.A1(\top.cb_syn.char_index[2] ),
    .A2(_03042_),
    .B1(\top.cb_syn.char_index[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03159_));
 sky130_fd_sc_hd__a32o_1 _06289_ (.A1(net545),
    .A2(_03045_),
    .A3(_03159_),
    .B1(_02583_),
    .B2(\top.cb_syn.curr_index[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03160_));
 sky130_fd_sc_hd__a21bo_1 _06290_ (.A1(net461),
    .A2(_03160_),
    .B1_N(_03158_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03161_));
 sky130_fd_sc_hd__a221o_1 _06291_ (.A1(net458),
    .A2(_03147_),
    .B1(_03152_),
    .B2(_02607_),
    .C1(_03161_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03162_));
 sky130_fd_sc_hd__a31o_1 _06292_ (.A1(net454),
    .A2(_03149_),
    .A3(_03151_),
    .B1(_03162_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03163_));
 sky130_fd_sc_hd__a22o_1 _06293_ (.A1(net1075),
    .A2(net165),
    .B1(_03163_),
    .B2(net208),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02127_));
 sky130_fd_sc_hd__or2_1 _06294_ (.A(net484),
    .B(_03089_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03164_));
 sky130_fd_sc_hd__a221o_1 _06295_ (.A1(net486),
    .A2(_02787_),
    .B1(_03090_),
    .B2(_03164_),
    .C1(_02601_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03165_));
 sky130_fd_sc_hd__xor2_1 _06296_ (.A(\top.cw1[4] ),
    .B(_03071_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03166_));
 sky130_fd_sc_hd__o211a_1 _06297_ (.A1(_02602_),
    .A2(_03166_),
    .B1(_03165_),
    .C1(net534),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03167_));
 sky130_fd_sc_hd__or3_1 _06298_ (.A(\top.cw2[4] ),
    .B(\top.cw2[3] ),
    .C(_03077_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03168_));
 sky130_fd_sc_hd__a32o_1 _06299_ (.A1(_02600_),
    .A2(_03079_),
    .A3(_03168_),
    .B1(net361),
    .B2(net486),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03169_));
 sky130_fd_sc_hd__o21a_1 _06300_ (.A1(_03167_),
    .A2(_03169_),
    .B1(net459),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03170_));
 sky130_fd_sc_hd__xnor2_1 _06301_ (.A(\top.sram_interface.init_counter[4] ),
    .B(_03020_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03171_));
 sky130_fd_sc_hd__xor2_1 _06302_ (.A(\top.hist_addr[4] ),
    .B(_03098_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03172_));
 sky130_fd_sc_hd__o221a_1 _06303_ (.A1(_03019_),
    .A2(_03171_),
    .B1(_03172_),
    .B2(\top.histogram.init ),
    .C1(net454),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03173_));
 sky130_fd_sc_hd__o22a_1 _06304_ (.A1(\top.cb_syn.char_index[2] ),
    .A2(\top.cb_syn.char_index[1] ),
    .B1(_02588_),
    .B2(net309),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03174_));
 sky130_fd_sc_hd__a22o_1 _06305_ (.A1(net545),
    .A2(_03043_),
    .B1(_03174_),
    .B2(_03034_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03175_));
 sky130_fd_sc_hd__o211a_1 _06306_ (.A1(\top.cb_syn.char_index[2] ),
    .A2(_03042_),
    .B1(_03175_),
    .C1(net465),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03176_));
 sky130_fd_sc_hd__or2_1 _06307_ (.A(net445),
    .B(\top.TRN_char_index[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03177_));
 sky130_fd_sc_hd__a32o_1 _06308_ (.A1(_02589_),
    .A2(_03049_),
    .A3(_03177_),
    .B1(_03054_),
    .B2(net545),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03178_));
 sky130_fd_sc_hd__o211a_1 _06309_ (.A1(net445),
    .A2(_03053_),
    .B1(_03178_),
    .C1(\top.controller.state_reg[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03179_));
 sky130_fd_sc_hd__a22o_1 _06310_ (.A1(\top.cb_syn.max_index[4] ),
    .A2(_03102_),
    .B1(_03104_),
    .B2(\top.hTree.nullSumIndex[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03180_));
 sky130_fd_sc_hd__a221o_1 _06311_ (.A1(\top.cb_syn.curr_index[4] ),
    .A2(_02584_),
    .B1(_03180_),
    .B2(net446),
    .C1(_03179_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03181_));
 sky130_fd_sc_hd__or4_1 _06312_ (.A(_03170_),
    .B(_03173_),
    .C(_03176_),
    .D(_03181_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03182_));
 sky130_fd_sc_hd__a22o_1 _06313_ (.A1(net68),
    .A2(net165),
    .B1(_03182_),
    .B2(net208),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02126_));
 sky130_fd_sc_hd__nand2_1 _06314_ (.A(\top.cw1[3] ),
    .B(_03070_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03183_));
 sky130_fd_sc_hd__nand2_1 _06315_ (.A(_03071_),
    .B(_03183_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03184_));
 sky130_fd_sc_hd__nand2_1 _06316_ (.A(net486),
    .B(_03088_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03185_));
 sky130_fd_sc_hd__nand3_1 _06317_ (.A(net406),
    .B(_03089_),
    .C(_03185_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03186_));
 sky130_fd_sc_hd__o211a_1 _06318_ (.A1(\top.findLeastValue.histo_index[2] ),
    .A2(net406),
    .B1(_03186_),
    .C1(net535),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03187_));
 sky130_fd_sc_hd__xnor2_1 _06319_ (.A(\top.cw2[3] ),
    .B(_03077_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03188_));
 sky130_fd_sc_hd__a221o_1 _06320_ (.A1(\top.findLeastValue.histo_index[2] ),
    .A2(net361),
    .B1(_02600_),
    .B2(_03188_),
    .C1(_03187_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03189_));
 sky130_fd_sc_hd__a21o_1 _06321_ (.A1(_02603_),
    .A2(_03184_),
    .B1(_03189_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03190_));
 sky130_fd_sc_hd__a22o_1 _06322_ (.A1(\top.cb_syn.max_index[3] ),
    .A2(_03102_),
    .B1(_03104_),
    .B2(\top.hTree.nullSumIndex[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03191_));
 sky130_fd_sc_hd__nand2_1 _06323_ (.A(\top.cb_syn.char_index[1] ),
    .B(\top.cb_syn.char_index[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03192_));
 sky130_fd_sc_hd__a21oi_1 _06324_ (.A1(_03042_),
    .A2(_03192_),
    .B1(_02605_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03193_));
 sky130_fd_sc_hd__nand2_1 _06325_ (.A(\top.TRN_char_index[1] ),
    .B(\top.TRN_char_index[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03194_));
 sky130_fd_sc_hd__a21oi_1 _06326_ (.A1(_03053_),
    .A2(_03194_),
    .B1(_02585_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03195_));
 sky130_fd_sc_hd__a2bb2o_1 _06327_ (.A1_N(\top.TRN_char_index[1] ),
    .A2_N(_02591_),
    .B1(_03191_),
    .B2(net446),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03196_));
 sky130_fd_sc_hd__or3_1 _06328_ (.A(_03193_),
    .B(_03195_),
    .C(_03196_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03197_));
 sky130_fd_sc_hd__a221o_1 _06329_ (.A1(\top.cb_syn.curr_index[3] ),
    .A2(_02584_),
    .B1(_02607_),
    .B2(_02537_),
    .C1(_03197_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03198_));
 sky130_fd_sc_hd__nand2_1 _06330_ (.A(_02416_),
    .B(_03098_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03199_));
 sky130_fd_sc_hd__a41o_1 _06331_ (.A1(\top.hist_addr[3] ),
    .A2(\top.hist_addr[2] ),
    .A3(\top.hist_addr[1] ),
    .A4(\top.hist_addr[0] ),
    .B1(_03199_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03200_));
 sky130_fd_sc_hd__o311a_1 _06332_ (.A1(_02927_),
    .A2(_03019_),
    .A3(_03020_),
    .B1(_03200_),
    .C1(net454),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03201_));
 sky130_fd_sc_hd__a211o_1 _06333_ (.A1(net458),
    .A2(_03190_),
    .B1(_03198_),
    .C1(_03201_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03202_));
 sky130_fd_sc_hd__a22o_1 _06334_ (.A1(net1077),
    .A2(net165),
    .B1(_03202_),
    .B2(net208),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02125_));
 sky130_fd_sc_hd__and2_1 _06335_ (.A(net487),
    .B(_02787_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03203_));
 sky130_fd_sc_hd__a21oi_1 _06336_ (.A1(net487),
    .A2(\top.findLeastValue.histo_index[0] ),
    .B1(\top.findLeastValue.histo_index[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03204_));
 sky130_fd_sc_hd__nor2_1 _06337_ (.A(_03088_),
    .B(_03204_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03205_));
 sky130_fd_sc_hd__a211o_1 _06338_ (.A1(net407),
    .A2(_03205_),
    .B1(_03203_),
    .C1(_02601_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03206_));
 sky130_fd_sc_hd__a21oi_1 _06339_ (.A1(\top.cw1[1] ),
    .A2(\top.cw1[0] ),
    .B1(\top.cw1[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03207_));
 sky130_fd_sc_hd__o21ai_1 _06340_ (.A1(_03070_),
    .A2(_03207_),
    .B1(_02601_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03208_));
 sky130_fd_sc_hd__nand2_1 _06341_ (.A(_02510_),
    .B(_03076_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03209_));
 sky130_fd_sc_hd__a32o_1 _06342_ (.A1(_02600_),
    .A2(_03078_),
    .A3(_03209_),
    .B1(_02578_),
    .B2(net487),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03210_));
 sky130_fd_sc_hd__a31o_1 _06343_ (.A1(net534),
    .A2(_03206_),
    .A3(_03208_),
    .B1(_03210_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03211_));
 sky130_fd_sc_hd__a21oi_1 _06344_ (.A1(\top.sram_interface.init_counter[1] ),
    .A2(\top.sram_interface.init_counter[0] ),
    .B1(\top.sram_interface.init_counter[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03212_));
 sky130_fd_sc_hd__nor2_1 _06345_ (.A(_02926_),
    .B(_03212_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03213_));
 sky130_fd_sc_hd__xnor2_1 _06346_ (.A(\top.hist_addr[2] ),
    .B(_03097_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03214_));
 sky130_fd_sc_hd__o221a_1 _06347_ (.A1(_03019_),
    .A2(_03213_),
    .B1(_03214_),
    .B2(\top.histogram.init ),
    .C1(net454),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03215_));
 sky130_fd_sc_hd__a22o_1 _06348_ (.A1(\top.cb_syn.max_index[2] ),
    .A2(_03102_),
    .B1(_03104_),
    .B2(\top.hTree.nullSumIndex[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03216_));
 sky130_fd_sc_hd__mux2_1 _06349_ (.A0(net545),
    .A1(_02589_),
    .S(\top.TRN_char_index[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03217_));
 sky130_fd_sc_hd__a2bb2o_1 _06350_ (.A1_N(\top.cb_syn.char_index[0] ),
    .A2_N(_02605_),
    .B1(_03217_),
    .B2(\top.controller.state_reg[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03218_));
 sky130_fd_sc_hd__a221o_1 _06351_ (.A1(\top.cb_syn.curr_index[2] ),
    .A2(_02584_),
    .B1(_03216_),
    .B2(net446),
    .C1(_03218_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03219_));
 sky130_fd_sc_hd__a21o_1 _06352_ (.A1(\top.cb_syn.char_index[0] ),
    .A2(_02607_),
    .B1(_03219_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03220_));
 sky130_fd_sc_hd__a211o_1 _06353_ (.A1(net458),
    .A2(_03211_),
    .B1(_03215_),
    .C1(_03220_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03221_));
 sky130_fd_sc_hd__a22o_1 _06354_ (.A1(net1261),
    .A2(net165),
    .B1(_03221_),
    .B2(net208),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02124_));
 sky130_fd_sc_hd__nand2_1 _06355_ (.A(_02574_),
    .B(_03087_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03222_));
 sky130_fd_sc_hd__o221ai_1 _06356_ (.A1(net406),
    .A2(_03087_),
    .B1(_03203_),
    .B2(_03222_),
    .C1(_02602_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03223_));
 sky130_fd_sc_hd__xor2_1 _06357_ (.A(\top.cw1[1] ),
    .B(\top.cw1[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03224_));
 sky130_fd_sc_hd__o211a_1 _06358_ (.A1(_02602_),
    .A2(_03224_),
    .B1(_03223_),
    .C1(net535),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03225_));
 sky130_fd_sc_hd__or2_1 _06359_ (.A(\top.cw2[1] ),
    .B(\top.cw2[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03226_));
 sky130_fd_sc_hd__a32o_1 _06360_ (.A1(_02600_),
    .A2(_03076_),
    .A3(_03226_),
    .B1(_02578_),
    .B2(\top.findLeastValue.histo_index[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03227_));
 sky130_fd_sc_hd__o21a_1 _06361_ (.A1(_03225_),
    .A2(_03227_),
    .B1(net459),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03228_));
 sky130_fd_sc_hd__xor2_1 _06362_ (.A(\top.sram_interface.init_counter[1] ),
    .B(\top.sram_interface.init_counter[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03229_));
 sky130_fd_sc_hd__or2_1 _06363_ (.A(\top.hist_addr[1] ),
    .B(\top.hist_addr[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03230_));
 sky130_fd_sc_hd__a21o_1 _06364_ (.A1(_03097_),
    .A2(_03230_),
    .B1(\top.histogram.init ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03231_));
 sky130_fd_sc_hd__o211a_1 _06365_ (.A1(_03019_),
    .A2(_03229_),
    .B1(_03231_),
    .C1(\top.controller.state_reg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03232_));
 sky130_fd_sc_hd__a22o_1 _06366_ (.A1(\top.cb_syn.max_index[1] ),
    .A2(_03102_),
    .B1(_03104_),
    .B2(\top.hTree.nullSumIndex[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03233_));
 sky130_fd_sc_hd__a221o_1 _06367_ (.A1(_02588_),
    .A2(_03013_),
    .B1(_03233_),
    .B2(net446),
    .C1(_03228_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03234_));
 sky130_fd_sc_hd__a211o_1 _06368_ (.A1(\top.cb_syn.curr_index[1] ),
    .A2(_02584_),
    .B1(_03232_),
    .C1(_03234_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03235_));
 sky130_fd_sc_hd__a22o_1 _06369_ (.A1(net1204),
    .A2(net165),
    .B1(_03235_),
    .B2(net208),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02123_));
 sky130_fd_sc_hd__a31o_1 _06370_ (.A1(_02504_),
    .A2(net534),
    .A3(net407),
    .B1(_02578_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03236_));
 sky130_fd_sc_hd__a221o_1 _06371_ (.A1(_02512_),
    .A2(_02600_),
    .B1(_02603_),
    .B2(_02513_),
    .C1(_03236_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03237_));
 sky130_fd_sc_hd__nand2_1 _06372_ (.A(net459),
    .B(_03237_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03238_));
 sky130_fd_sc_hd__a221o_1 _06373_ (.A1(_02416_),
    .A2(\top.hist_addr[0] ),
    .B1(_03018_),
    .B2(\top.sram_interface.init_counter[0] ),
    .C1(_02417_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03239_));
 sky130_fd_sc_hd__o21a_1 _06374_ (.A1(net528),
    .A2(net309),
    .B1(net461),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03240_));
 sky130_fd_sc_hd__a221o_1 _06375_ (.A1(net460),
    .A2(\top.sram_interface.word_cnt[9] ),
    .B1(_02586_),
    .B2(net451),
    .C1(_02862_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03241_));
 sky130_fd_sc_hd__or4bb_1 _06376_ (.A(_03241_),
    .B(_03240_),
    .C_N(_03239_),
    .D_N(_03238_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03242_));
 sky130_fd_sc_hd__a22o_1 _06377_ (.A1(net1174),
    .A2(net164),
    .B1(_03242_),
    .B2(net208),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02122_));
 sky130_fd_sc_hd__and3_4 _06378_ (.A(net439),
    .B(\top.histogram.state[3] ),
    .C(net360),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03243_));
 sky130_fd_sc_hd__or3b_4 _06379_ (.A(_02594_),
    .B(net444),
    .C_N(\top.histogram.state[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03244_));
 sky130_fd_sc_hd__nand2_1 _06380_ (.A(\top.hist_data_o[1] ),
    .B(\top.hist_data_o[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03245_));
 sky130_fd_sc_hd__and4_1 _06381_ (.A(\top.hist_data_o[3] ),
    .B(\top.hist_data_o[2] ),
    .C(\top.hist_data_o[1] ),
    .D(\top.hist_data_o[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03246_));
 sky130_fd_sc_hd__and2_1 _06382_ (.A(\top.hist_data_o[5] ),
    .B(\top.hist_data_o[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03247_));
 sky130_fd_sc_hd__and2_1 _06383_ (.A(_03246_),
    .B(_03247_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03248_));
 sky130_fd_sc_hd__and3_2 _06384_ (.A(\top.hist_data_o[7] ),
    .B(\top.hist_data_o[6] ),
    .C(_03248_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03249_));
 sky130_fd_sc_hd__and2_1 _06385_ (.A(\top.hist_data_o[8] ),
    .B(_03249_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03250_));
 sky130_fd_sc_hd__and3_1 _06386_ (.A(\top.hist_data_o[10] ),
    .B(\top.hist_data_o[9] ),
    .C(_03250_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03251_));
 sky130_fd_sc_hd__and4_1 _06387_ (.A(\top.hist_data_o[11] ),
    .B(\top.hist_data_o[10] ),
    .C(\top.hist_data_o[9] ),
    .D(\top.hist_data_o[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03252_));
 sky130_fd_sc_hd__and3_1 _06388_ (.A(\top.hist_data_o[12] ),
    .B(_03249_),
    .C(_03252_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03253_));
 sky130_fd_sc_hd__and2_1 _06389_ (.A(\top.hist_data_o[13] ),
    .B(\top.hist_data_o[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03254_));
 sky130_fd_sc_hd__and3_1 _06390_ (.A(_03249_),
    .B(_03252_),
    .C(_03254_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03255_));
 sky130_fd_sc_hd__and4_1 _06391_ (.A(\top.hist_data_o[14] ),
    .B(_03249_),
    .C(_03252_),
    .D(_03254_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03256_));
 sky130_fd_sc_hd__and4_1 _06392_ (.A(\top.hist_data_o[17] ),
    .B(\top.hist_data_o[16] ),
    .C(\top.hist_data_o[15] ),
    .D(_03256_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03257_));
 sky130_fd_sc_hd__and4_1 _06393_ (.A(\top.hist_data_o[20] ),
    .B(\top.hist_data_o[19] ),
    .C(\top.hist_data_o[18] ),
    .D(_03257_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03258_));
 sky130_fd_sc_hd__and3_1 _06394_ (.A(\top.hist_data_o[22] ),
    .B(\top.hist_data_o[21] ),
    .C(_03258_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03259_));
 sky130_fd_sc_hd__and2_1 _06395_ (.A(\top.hist_data_o[23] ),
    .B(_03259_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03260_));
 sky130_fd_sc_hd__and3_1 _06396_ (.A(\top.hist_data_o[25] ),
    .B(\top.hist_data_o[24] ),
    .C(_03260_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03261_));
 sky130_fd_sc_hd__and2_1 _06397_ (.A(\top.hist_data_o[26] ),
    .B(_03261_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03262_));
 sky130_fd_sc_hd__and3_1 _06398_ (.A(\top.hist_data_o[28] ),
    .B(\top.hist_data_o[27] ),
    .C(_03262_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03263_));
 sky130_fd_sc_hd__and2_1 _06399_ (.A(\top.hist_data_o[29] ),
    .B(_03263_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03264_));
 sky130_fd_sc_hd__nand2_1 _06400_ (.A(\top.hist_data_o[30] ),
    .B(_03264_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03265_));
 sky130_fd_sc_hd__and3_1 _06401_ (.A(\top.hist_data_o[15] ),
    .B(\top.hist_data_o[14] ),
    .C(_03255_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03266_));
 sky130_fd_sc_hd__and2_1 _06402_ (.A(\top.hist_data_o[16] ),
    .B(_03266_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03267_));
 sky130_fd_sc_hd__and3_1 _06403_ (.A(\top.hist_data_o[18] ),
    .B(\top.hist_data_o[17] ),
    .C(_03267_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03268_));
 sky130_fd_sc_hd__and3_1 _06404_ (.A(\top.hist_data_o[20] ),
    .B(\top.hist_data_o[19] ),
    .C(_03268_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03269_));
 sky130_fd_sc_hd__xnor2_1 _06405_ (.A(\top.hist_data_o[31] ),
    .B(_03265_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03270_));
 sky130_fd_sc_hd__mux2_1 _06406_ (.A0(net1429),
    .A1(_03270_),
    .S(net301),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02121_));
 sky130_fd_sc_hd__and3_1 _06407_ (.A(\top.hist_data_o[17] ),
    .B(\top.hist_data_o[16] ),
    .C(_03266_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03271_));
 sky130_fd_sc_hd__and3_1 _06408_ (.A(\top.hist_data_o[19] ),
    .B(\top.hist_data_o[18] ),
    .C(_03271_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03272_));
 sky130_fd_sc_hd__and3_1 _06409_ (.A(\top.hist_data_o[21] ),
    .B(\top.hist_data_o[20] ),
    .C(_03272_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03273_));
 sky130_fd_sc_hd__xor2_1 _06410_ (.A(\top.hist_data_o[30] ),
    .B(_03264_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03274_));
 sky130_fd_sc_hd__mux2_1 _06411_ (.A0(net1251),
    .A1(_03274_),
    .S(net301),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02120_));
 sky130_fd_sc_hd__nor2_1 _06412_ (.A(\top.hist_data_o[29] ),
    .B(_03263_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03275_));
 sky130_fd_sc_hd__o21ai_1 _06413_ (.A1(_03264_),
    .A2(_03275_),
    .B1(net301),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03276_));
 sky130_fd_sc_hd__o21a_1 _06414_ (.A1(net1461),
    .A2(net301),
    .B1(_03276_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02119_));
 sky130_fd_sc_hd__a21oi_1 _06415_ (.A1(\top.hist_data_o[27] ),
    .A2(_03262_),
    .B1(\top.hist_data_o[28] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03277_));
 sky130_fd_sc_hd__nor2_1 _06416_ (.A(_03263_),
    .B(_03277_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03278_));
 sky130_fd_sc_hd__mux2_1 _06417_ (.A0(net1118),
    .A1(_03278_),
    .S(net301),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02118_));
 sky130_fd_sc_hd__xor2_1 _06418_ (.A(\top.hist_data_o[27] ),
    .B(_03262_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03279_));
 sky130_fd_sc_hd__mux2_1 _06419_ (.A0(net1653),
    .A1(_03279_),
    .S(net301),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02117_));
 sky130_fd_sc_hd__nor2_1 _06420_ (.A(\top.hist_data_o[26] ),
    .B(_03261_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03280_));
 sky130_fd_sc_hd__nor2_1 _06421_ (.A(_03262_),
    .B(_03280_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03281_));
 sky130_fd_sc_hd__mux2_1 _06422_ (.A0(net1180),
    .A1(_03281_),
    .S(net301),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02116_));
 sky130_fd_sc_hd__a21oi_1 _06423_ (.A1(\top.hist_data_o[24] ),
    .A2(_03260_),
    .B1(\top.hist_data_o[25] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03282_));
 sky130_fd_sc_hd__nor2_1 _06424_ (.A(_03261_),
    .B(_03282_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03283_));
 sky130_fd_sc_hd__mux2_1 _06425_ (.A0(net1126),
    .A1(_03283_),
    .S(net301),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02115_));
 sky130_fd_sc_hd__xor2_1 _06426_ (.A(\top.hist_data_o[24] ),
    .B(_03260_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03284_));
 sky130_fd_sc_hd__mux2_1 _06427_ (.A0(net1353),
    .A1(_03284_),
    .S(net301),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02114_));
 sky130_fd_sc_hd__or2_1 _06428_ (.A(\top.hist_data_o[23] ),
    .B(_03259_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03285_));
 sky130_fd_sc_hd__and3b_1 _06429_ (.A_N(_03260_),
    .B(_03285_),
    .C(net301),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03286_));
 sky130_fd_sc_hd__a21o_1 _06430_ (.A1(net1045),
    .A2(net299),
    .B1(_03286_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02113_));
 sky130_fd_sc_hd__o21ba_1 _06431_ (.A1(\top.hist_data_o[22] ),
    .A2(_03273_),
    .B1_N(_03259_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03287_));
 sky130_fd_sc_hd__mux2_1 _06432_ (.A0(net1188),
    .A1(_03287_),
    .S(net300),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02112_));
 sky130_fd_sc_hd__o21ba_1 _06433_ (.A1(\top.hist_data_o[21] ),
    .A2(_03269_),
    .B1_N(_03273_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03288_));
 sky130_fd_sc_hd__mux2_1 _06434_ (.A0(net1145),
    .A1(_03288_),
    .S(_03243_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02111_));
 sky130_fd_sc_hd__o21ba_1 _06435_ (.A1(\top.hist_data_o[20] ),
    .A2(_03272_),
    .B1_N(_03258_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03289_));
 sky130_fd_sc_hd__mux2_1 _06436_ (.A0(net1167),
    .A1(_03289_),
    .S(net300),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02110_));
 sky130_fd_sc_hd__o21ba_1 _06437_ (.A1(\top.hist_data_o[19] ),
    .A2(_03268_),
    .B1_N(_03272_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03290_));
 sky130_fd_sc_hd__mux2_1 _06438_ (.A0(net1108),
    .A1(_03290_),
    .S(net300),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02109_));
 sky130_fd_sc_hd__o21ba_1 _06439_ (.A1(\top.hist_data_o[18] ),
    .A2(_03271_),
    .B1_N(_03268_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03291_));
 sky130_fd_sc_hd__mux2_1 _06440_ (.A0(net1140),
    .A1(_03291_),
    .S(net300),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02108_));
 sky130_fd_sc_hd__o21ba_1 _06441_ (.A1(\top.hist_data_o[17] ),
    .A2(_03267_),
    .B1_N(_03271_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03292_));
 sky130_fd_sc_hd__mux2_1 _06442_ (.A0(net1305),
    .A1(_03292_),
    .S(_03243_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02107_));
 sky130_fd_sc_hd__nor2_1 _06443_ (.A(\top.hist_data_o[16] ),
    .B(_03266_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03293_));
 sky130_fd_sc_hd__nand2_1 _06444_ (.A(net1058),
    .B(net298),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03294_));
 sky130_fd_sc_hd__o31ai_1 _06445_ (.A1(net298),
    .A2(_03267_),
    .A3(_03293_),
    .B1(_03294_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02106_));
 sky130_fd_sc_hd__xor2_1 _06446_ (.A(\top.hist_data_o[15] ),
    .B(_03256_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03295_));
 sky130_fd_sc_hd__mux2_1 _06447_ (.A0(net1125),
    .A1(_03295_),
    .S(net300),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02105_));
 sky130_fd_sc_hd__nor2_1 _06448_ (.A(\top.hist_data_o[14] ),
    .B(_03255_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03296_));
 sky130_fd_sc_hd__nand2_1 _06449_ (.A(net1013),
    .B(net298),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03297_));
 sky130_fd_sc_hd__o31ai_1 _06450_ (.A1(net298),
    .A2(_03256_),
    .A3(_03296_),
    .B1(_03297_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02104_));
 sky130_fd_sc_hd__nor2_1 _06451_ (.A(\top.hist_data_o[13] ),
    .B(_03253_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03298_));
 sky130_fd_sc_hd__nand2_1 _06452_ (.A(net1312),
    .B(net298),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03299_));
 sky130_fd_sc_hd__o31ai_1 _06453_ (.A1(net298),
    .A2(_03255_),
    .A3(_03298_),
    .B1(_03299_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02103_));
 sky130_fd_sc_hd__a21oi_1 _06454_ (.A1(_03249_),
    .A2(_03252_),
    .B1(\top.hist_data_o[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03300_));
 sky130_fd_sc_hd__nand2_1 _06455_ (.A(net1472),
    .B(net298),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03301_));
 sky130_fd_sc_hd__o31ai_1 _06456_ (.A1(net299),
    .A2(_03253_),
    .A3(_03300_),
    .B1(_03301_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02102_));
 sky130_fd_sc_hd__nor2_1 _06457_ (.A(\top.hist_data_o[11] ),
    .B(_03251_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03302_));
 sky130_fd_sc_hd__a21oi_1 _06458_ (.A1(_03249_),
    .A2(_03252_),
    .B1(_03302_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03303_));
 sky130_fd_sc_hd__mux2_1 _06459_ (.A0(net1366),
    .A1(_03303_),
    .S(net300),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02101_));
 sky130_fd_sc_hd__a31o_1 _06460_ (.A1(\top.hist_data_o[9] ),
    .A2(\top.hist_data_o[8] ),
    .A3(_03249_),
    .B1(\top.hist_data_o[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03304_));
 sky130_fd_sc_hd__nor2_1 _06461_ (.A(net299),
    .B(_03251_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03305_));
 sky130_fd_sc_hd__a22o_1 _06462_ (.A1(net1576),
    .A2(net299),
    .B1(_03304_),
    .B2(_03305_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02100_));
 sky130_fd_sc_hd__xor2_1 _06463_ (.A(\top.hist_data_o[9] ),
    .B(_03250_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03306_));
 sky130_fd_sc_hd__mux2_1 _06464_ (.A0(net1278),
    .A1(_03306_),
    .S(net300),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02099_));
 sky130_fd_sc_hd__nor2_1 _06465_ (.A(\top.hist_data_o[8] ),
    .B(_03249_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03307_));
 sky130_fd_sc_hd__nor2_1 _06466_ (.A(_03250_),
    .B(_03307_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03308_));
 sky130_fd_sc_hd__mux2_1 _06467_ (.A0(net1467),
    .A1(_03308_),
    .S(net300),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02098_));
 sky130_fd_sc_hd__a31o_1 _06468_ (.A1(\top.hist_data_o[6] ),
    .A2(_03246_),
    .A3(_03247_),
    .B1(\top.hist_data_o[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03309_));
 sky130_fd_sc_hd__nor2_1 _06469_ (.A(net298),
    .B(_03249_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03310_));
 sky130_fd_sc_hd__a22o_1 _06470_ (.A1(net1527),
    .A2(net297),
    .B1(_03309_),
    .B2(_03310_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02097_));
 sky130_fd_sc_hd__a21oi_1 _06471_ (.A1(\top.hist_data_o[6] ),
    .A2(_03248_),
    .B1(net298),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03311_));
 sky130_fd_sc_hd__o21a_1 _06472_ (.A1(\top.hist_data_o[6] ),
    .A2(_03248_),
    .B1(_03311_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03312_));
 sky130_fd_sc_hd__a21o_1 _06473_ (.A1(net1376),
    .A2(net297),
    .B1(_03312_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02096_));
 sky130_fd_sc_hd__a21o_1 _06474_ (.A1(\top.hist_data_o[4] ),
    .A2(_03246_),
    .B1(\top.hist_data_o[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03313_));
 sky130_fd_sc_hd__nor2_1 _06475_ (.A(net297),
    .B(_03248_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03314_));
 sky130_fd_sc_hd__a22o_1 _06476_ (.A1(net1464),
    .A2(net297),
    .B1(_03313_),
    .B2(_03314_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02095_));
 sky130_fd_sc_hd__a21oi_1 _06477_ (.A1(\top.hist_data_o[4] ),
    .A2(_03246_),
    .B1(net297),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03315_));
 sky130_fd_sc_hd__o21a_1 _06478_ (.A1(\top.hist_data_o[4] ),
    .A2(_03246_),
    .B1(_03315_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03316_));
 sky130_fd_sc_hd__a21o_1 _06479_ (.A1(net1155),
    .A2(net297),
    .B1(_03316_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02094_));
 sky130_fd_sc_hd__a31o_1 _06480_ (.A1(\top.hist_data_o[2] ),
    .A2(\top.hist_data_o[1] ),
    .A3(\top.hist_data_o[0] ),
    .B1(\top.hist_data_o[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03317_));
 sky130_fd_sc_hd__nor2_1 _06481_ (.A(net297),
    .B(_03246_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03318_));
 sky130_fd_sc_hd__a22o_1 _06482_ (.A1(net1346),
    .A2(net297),
    .B1(_03317_),
    .B2(_03318_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02093_));
 sky130_fd_sc_hd__xnor2_1 _06483_ (.A(\top.hist_data_o[2] ),
    .B(_03245_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03319_));
 sky130_fd_sc_hd__mux2_1 _06484_ (.A0(net1498),
    .A1(_03319_),
    .S(net300),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02092_));
 sky130_fd_sc_hd__o21a_1 _06485_ (.A1(\top.hist_data_o[1] ),
    .A2(\top.hist_data_o[0] ),
    .B1(net300),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03320_));
 sky130_fd_sc_hd__a22o_1 _06486_ (.A1(net1410),
    .A2(net297),
    .B1(_03245_),
    .B2(_03320_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02091_));
 sky130_fd_sc_hd__mux2_1 _06487_ (.A0(_02420_),
    .A1(net1454),
    .S(net297),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02090_));
 sky130_fd_sc_hd__and2b_1 _06488_ (.A_N(\top.dut.out_valid ),
    .B(\top.histogram.out_of_init ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03321_));
 sky130_fd_sc_hd__or2_1 _06489_ (.A(_02454_),
    .B(_03321_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03322_));
 sky130_fd_sc_hd__o21a_1 _06490_ (.A1(\top.histogram.eof_n ),
    .A2(\top.histogram.state[1] ),
    .B1(net453),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03323_));
 sky130_fd_sc_hd__and2_1 _06491_ (.A(_03322_),
    .B(_03323_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03324_));
 sky130_fd_sc_hd__o2111a_2 _06492_ (.A1(_02454_),
    .A2(_03321_),
    .B1(_03323_),
    .C1(\top.histogram.total[0] ),
    .D1(\top.histogram.total[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03325_));
 sky130_fd_sc_hd__and3_1 _06493_ (.A(\top.histogram.total[3] ),
    .B(\top.histogram.total[2] ),
    .C(_03325_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03326_));
 sky130_fd_sc_hd__and2_1 _06494_ (.A(\top.histogram.total[4] ),
    .B(_03326_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03327_));
 sky130_fd_sc_hd__and4_1 _06495_ (.A(\top.histogram.total[5] ),
    .B(\top.histogram.total[4] ),
    .C(\top.histogram.total[3] ),
    .D(\top.histogram.total[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03328_));
 sky130_fd_sc_hd__and3_1 _06496_ (.A(\top.histogram.total[6] ),
    .B(_03325_),
    .C(_03328_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03329_));
 sky130_fd_sc_hd__and2_1 _06497_ (.A(\top.histogram.total[7] ),
    .B(\top.histogram.total[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03330_));
 sky130_fd_sc_hd__and4_1 _06498_ (.A(\top.histogram.total[8] ),
    .B(_03325_),
    .C(_03328_),
    .D(_03330_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03331_));
 sky130_fd_sc_hd__and4_1 _06499_ (.A(\top.histogram.total[11] ),
    .B(\top.histogram.total[10] ),
    .C(\top.histogram.total[9] ),
    .D(_03331_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03332_));
 sky130_fd_sc_hd__and3_1 _06500_ (.A(\top.histogram.total[13] ),
    .B(\top.histogram.total[12] ),
    .C(_03332_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03333_));
 sky130_fd_sc_hd__and4_1 _06501_ (.A(\top.histogram.total[16] ),
    .B(\top.histogram.total[15] ),
    .C(\top.histogram.total[14] ),
    .D(_03333_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03334_));
 sky130_fd_sc_hd__and3_1 _06502_ (.A(\top.histogram.total[18] ),
    .B(\top.histogram.total[17] ),
    .C(_03334_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03335_));
 sky130_fd_sc_hd__and3_1 _06503_ (.A(\top.histogram.total[20] ),
    .B(\top.histogram.total[19] ),
    .C(_03335_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03336_));
 sky130_fd_sc_hd__and2_1 _06504_ (.A(\top.histogram.total[21] ),
    .B(_03336_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03337_));
 sky130_fd_sc_hd__and3_1 _06505_ (.A(\top.histogram.total[22] ),
    .B(\top.histogram.total[21] ),
    .C(_03336_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03338_));
 sky130_fd_sc_hd__and3_1 _06506_ (.A(\top.histogram.total[24] ),
    .B(\top.histogram.total[23] ),
    .C(_03338_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03339_));
 sky130_fd_sc_hd__and2_1 _06507_ (.A(\top.histogram.total[25] ),
    .B(_03339_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03340_));
 sky130_fd_sc_hd__and3_1 _06508_ (.A(\top.histogram.total[27] ),
    .B(\top.histogram.total[26] ),
    .C(_03340_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03341_));
 sky130_fd_sc_hd__and3_1 _06509_ (.A(\top.histogram.total[29] ),
    .B(\top.histogram.total[28] ),
    .C(_03341_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03342_));
 sky130_fd_sc_hd__nand2_1 _06510_ (.A(\top.histogram.total[30] ),
    .B(_03342_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03343_));
 sky130_fd_sc_hd__and3b_1 _06511_ (.A_N(\top.histogram.total[31] ),
    .B(\top.histogram.total[30] ),
    .C(_03342_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03344_));
 sky130_fd_sc_hd__a21o_1 _06512_ (.A1(net1364),
    .A2(_03343_),
    .B1(_03344_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02089_));
 sky130_fd_sc_hd__xor2_1 _06513_ (.A(net1501),
    .B(_03342_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02088_));
 sky130_fd_sc_hd__a21oi_1 _06514_ (.A1(\top.histogram.total[28] ),
    .A2(_03341_),
    .B1(net1448),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03345_));
 sky130_fd_sc_hd__nor2_1 _06515_ (.A(_03342_),
    .B(net1449),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02087_));
 sky130_fd_sc_hd__xor2_1 _06516_ (.A(net1505),
    .B(_03341_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02086_));
 sky130_fd_sc_hd__a21oi_1 _06517_ (.A1(\top.histogram.total[26] ),
    .A2(_03340_),
    .B1(net1506),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03346_));
 sky130_fd_sc_hd__nor2_1 _06518_ (.A(_03341_),
    .B(net1507),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02085_));
 sky130_fd_sc_hd__xor2_1 _06519_ (.A(net1487),
    .B(_03340_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02084_));
 sky130_fd_sc_hd__nor2_1 _06520_ (.A(net1611),
    .B(_03339_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03347_));
 sky130_fd_sc_hd__nor2_1 _06521_ (.A(_03340_),
    .B(_03347_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02083_));
 sky130_fd_sc_hd__a21oi_1 _06522_ (.A1(\top.histogram.total[23] ),
    .A2(_03338_),
    .B1(net1544),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03348_));
 sky130_fd_sc_hd__nor2_1 _06523_ (.A(_03339_),
    .B(net1545),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02082_));
 sky130_fd_sc_hd__xor2_1 _06524_ (.A(net1456),
    .B(_03338_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02081_));
 sky130_fd_sc_hd__nor2_1 _06525_ (.A(net1532),
    .B(_03337_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03349_));
 sky130_fd_sc_hd__nor2_1 _06526_ (.A(_03338_),
    .B(_03349_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02080_));
 sky130_fd_sc_hd__nor2_1 _06527_ (.A(net1643),
    .B(_03336_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03350_));
 sky130_fd_sc_hd__nor2_1 _06528_ (.A(_03337_),
    .B(_03350_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02079_));
 sky130_fd_sc_hd__a21oi_1 _06529_ (.A1(\top.histogram.total[19] ),
    .A2(_03335_),
    .B1(net1520),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03351_));
 sky130_fd_sc_hd__nor2_1 _06530_ (.A(_03336_),
    .B(net1521),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02078_));
 sky130_fd_sc_hd__xor2_1 _06531_ (.A(net1512),
    .B(_03335_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02077_));
 sky130_fd_sc_hd__a21oi_1 _06532_ (.A1(net1798),
    .A2(_03334_),
    .B1(net1502),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03352_));
 sky130_fd_sc_hd__nor2_1 _06533_ (.A(_03335_),
    .B(_03352_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02076_));
 sky130_fd_sc_hd__xor2_1 _06534_ (.A(net1563),
    .B(_03334_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02075_));
 sky130_fd_sc_hd__and3_1 _06535_ (.A(\top.histogram.total[15] ),
    .B(\top.histogram.total[14] ),
    .C(_03333_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03353_));
 sky130_fd_sc_hd__o21ba_1 _06536_ (.A1(net1596),
    .A2(_03353_),
    .B1_N(_03334_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02074_));
 sky130_fd_sc_hd__a21oi_1 _06537_ (.A1(net1803),
    .A2(_03333_),
    .B1(net1591),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03354_));
 sky130_fd_sc_hd__nor2_1 _06538_ (.A(_03353_),
    .B(_03354_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02073_));
 sky130_fd_sc_hd__xor2_1 _06539_ (.A(net1597),
    .B(_03333_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02072_));
 sky130_fd_sc_hd__a21oi_1 _06540_ (.A1(\top.histogram.total[12] ),
    .A2(_03332_),
    .B1(net1503),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03355_));
 sky130_fd_sc_hd__nor2_1 _06541_ (.A(_03333_),
    .B(net1504),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02071_));
 sky130_fd_sc_hd__xor2_1 _06542_ (.A(net1478),
    .B(_03332_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02070_));
 sky130_fd_sc_hd__and3_1 _06543_ (.A(\top.histogram.total[10] ),
    .B(\top.histogram.total[9] ),
    .C(_03331_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03356_));
 sky130_fd_sc_hd__o21ba_1 _06544_ (.A1(net1519),
    .A2(_03356_),
    .B1_N(_03332_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02069_));
 sky130_fd_sc_hd__a21oi_1 _06545_ (.A1(\top.histogram.total[9] ),
    .A2(_03331_),
    .B1(net1632),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03357_));
 sky130_fd_sc_hd__nor2_1 _06546_ (.A(_03356_),
    .B(_03357_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02068_));
 sky130_fd_sc_hd__xor2_1 _06547_ (.A(net1593),
    .B(_03331_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02067_));
 sky130_fd_sc_hd__a31o_1 _06548_ (.A1(_03325_),
    .A2(_03328_),
    .A3(_03330_),
    .B1(\top.histogram.total[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03358_));
 sky130_fd_sc_hd__and2b_1 _06549_ (.A_N(_03331_),
    .B(_03358_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02066_));
 sky130_fd_sc_hd__xor2_1 _06550_ (.A(net1105),
    .B(_03329_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02065_));
 sky130_fd_sc_hd__a21oi_1 _06551_ (.A1(_03325_),
    .A2(_03328_),
    .B1(net1583),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03359_));
 sky130_fd_sc_hd__nor2_1 _06552_ (.A(_03329_),
    .B(_03359_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02064_));
 sky130_fd_sc_hd__nor2_1 _06553_ (.A(net1422),
    .B(_03327_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03360_));
 sky130_fd_sc_hd__a21oi_1 _06554_ (.A1(_03325_),
    .A2(_03328_),
    .B1(_03360_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02063_));
 sky130_fd_sc_hd__nor2_1 _06555_ (.A(net1668),
    .B(_03326_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03361_));
 sky130_fd_sc_hd__nor2_1 _06556_ (.A(_03327_),
    .B(_03361_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02062_));
 sky130_fd_sc_hd__a21oi_1 _06557_ (.A1(\top.histogram.total[2] ),
    .A2(_03325_),
    .B1(net1608),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03362_));
 sky130_fd_sc_hd__nor2_1 _06558_ (.A(_03326_),
    .B(net1609),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02061_));
 sky130_fd_sc_hd__xor2_1 _06559_ (.A(net1602),
    .B(_03325_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02060_));
 sky130_fd_sc_hd__a31o_1 _06560_ (.A1(\top.histogram.total[0] ),
    .A2(_03322_),
    .A3(_03323_),
    .B1(\top.histogram.total[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03363_));
 sky130_fd_sc_hd__and2b_1 _06561_ (.A_N(_03325_),
    .B(_03363_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02059_));
 sky130_fd_sc_hd__xor2_1 _06562_ (.A(net1578),
    .B(_03324_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02058_));
 sky130_fd_sc_hd__and2_1 _06563_ (.A(_02454_),
    .B(\top.histogram.state[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03364_));
 sky130_fd_sc_hd__a21bo_1 _06564_ (.A1(net453),
    .A2(_03364_),
    .B1_N(\top.controller.fin_HG ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03365_));
 sky130_fd_sc_hd__or4b_1 _06565_ (.A(\top.dut.out[7] ),
    .B(\top.dut.out[6] ),
    .C(\top.dut.out[5] ),
    .D_N(\top.dut.out[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03366_));
 sky130_fd_sc_hd__nor2_1 _06566_ (.A(\top.dut.out[0] ),
    .B(_03366_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03367_));
 sky130_fd_sc_hd__and4b_1 _06567_ (.A_N(\top.dut.out[2] ),
    .B(\top.dut.out[1] ),
    .C(_03367_),
    .D(\top.dut.out[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03368_));
 sky130_fd_sc_hd__or4b_1 _06568_ (.A(_02417_),
    .B(_02454_),
    .C(_02561_),
    .D_N(_03368_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03369_));
 sky130_fd_sc_hd__nand2_1 _06569_ (.A(_03365_),
    .B(_03369_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02057_));
 sky130_fd_sc_hd__and2_1 _06570_ (.A(\top.header_synthesis.write_char_path ),
    .B(\top.header_synthesis.start ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03370_));
 sky130_fd_sc_hd__nand2_1 _06571_ (.A(\top.header_synthesis.write_char_path ),
    .B(\top.header_synthesis.start ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03371_));
 sky130_fd_sc_hd__and3_1 _06572_ (.A(\top.header_synthesis.enable ),
    .B(\top.header_synthesis.write_char_path ),
    .C(\top.header_synthesis.char_added ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03372_));
 sky130_fd_sc_hd__or4_1 _06573_ (.A(\top.header_synthesis.count[7] ),
    .B(\top.header_synthesis.count[6] ),
    .C(\top.header_synthesis.count[5] ),
    .D(\top.header_synthesis.count[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03373_));
 sky130_fd_sc_hd__or3_1 _06574_ (.A(\top.header_synthesis.count[2] ),
    .B(\top.header_synthesis.count[1] ),
    .C(\top.header_synthesis.count[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03374_));
 sky130_fd_sc_hd__a21oi_2 _06575_ (.A1(\top.header_synthesis.count[3] ),
    .A2(_03374_),
    .B1(_03373_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03375_));
 sky130_fd_sc_hd__a21oi_1 _06576_ (.A1(_03372_),
    .A2(_03375_),
    .B1(_03370_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03376_));
 sky130_fd_sc_hd__and2b_1 _06577_ (.A_N(net296),
    .B(\top.header_synthesis.header[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03377_));
 sky130_fd_sc_hd__mux4_1 _06578_ (.A0(\top.cb_syn.num_lefts[0] ),
    .A1(\top.cb_syn.num_lefts[4] ),
    .A2(\top.cb_syn.num_lefts[6] ),
    .A3(\top.cb_syn.num_lefts[2] ),
    .S0(\top.header_synthesis.count[2] ),
    .S1(\top.header_synthesis.count[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03378_));
 sky130_fd_sc_hd__or2_1 _06579_ (.A(\top.header_synthesis.count[0] ),
    .B(_03378_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03379_));
 sky130_fd_sc_hd__mux4_1 _06580_ (.A0(\top.cb_syn.num_lefts[7] ),
    .A1(\top.cb_syn.num_lefts[5] ),
    .A2(\top.cb_syn.num_lefts[3] ),
    .A3(\top.cb_syn.num_lefts[1] ),
    .S0(\top.header_synthesis.count[1] ),
    .S1(\top.header_synthesis.count[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03380_));
 sky130_fd_sc_hd__o211a_1 _06581_ (.A1(_02544_),
    .A2(_03380_),
    .B1(_03379_),
    .C1(_03375_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03381_));
 sky130_fd_sc_hd__or3_1 _06582_ (.A(\top.header_synthesis.count[3] ),
    .B(_03373_),
    .C(_03374_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03382_));
 sky130_fd_sc_hd__nand2_1 _06583_ (.A(\top.header_synthesis.write_num_lefts ),
    .B(_03382_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03383_));
 sky130_fd_sc_hd__o22a_1 _06584_ (.A1(\top.header_synthesis.write_num_lefts ),
    .A2(_03377_),
    .B1(_03381_),
    .B2(_03383_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03384_));
 sky130_fd_sc_hd__or4_1 _06585_ (.A(\top.cb_syn.zeroes[5] ),
    .B(\top.cb_syn.zeroes[4] ),
    .C(\top.cb_syn.zeroes[3] ),
    .D(\top.cb_syn.zeroes[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03385_));
 sky130_fd_sc_hd__or2_1 _06586_ (.A(\top.cb_syn.zeroes[1] ),
    .B(\top.cb_syn.zeroes[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03386_));
 sky130_fd_sc_hd__or4_1 _06587_ (.A(\top.cb_syn.zeroes[7] ),
    .B(\top.cb_syn.zeroes[6] ),
    .C(_03385_),
    .D(_03386_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03387_));
 sky130_fd_sc_hd__nand2_2 _06588_ (.A(\top.cb_syn.state8 ),
    .B(_03387_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03388_));
 sky130_fd_sc_hd__nor2_1 _06589_ (.A(\top.header_synthesis.write_num_lefts ),
    .B(\top.header_synthesis.write_char_path ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03389_));
 sky130_fd_sc_hd__a31o_1 _06590_ (.A1(\top.header_synthesis.bit1 ),
    .A2(_03388_),
    .A3(_03389_),
    .B1(_03384_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02056_));
 sky130_fd_sc_hd__nand2_1 _06591_ (.A(_02843_),
    .B(_02852_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03390_));
 sky130_fd_sc_hd__and3_1 _06592_ (.A(net448),
    .B(net544),
    .C(_03390_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03391_));
 sky130_fd_sc_hd__or3b_1 _06593_ (.A(net431),
    .B(_02553_),
    .C_N(_03390_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03392_));
 sky130_fd_sc_hd__nor2_2 _06594_ (.A(_02865_),
    .B(_03392_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03393_));
 sky130_fd_sc_hd__or2_2 _06595_ (.A(_02865_),
    .B(_03392_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03394_));
 sky130_fd_sc_hd__nor2_1 _06596_ (.A(_02562_),
    .B(net288),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03395_));
 sky130_fd_sc_hd__a21o_1 _06597_ (.A1(\top.findLeastValue.startup ),
    .A2(_02562_),
    .B1(net288),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02055_));
 sky130_fd_sc_hd__or4_1 _06598_ (.A(\top.compVal[11] ),
    .B(\top.compVal[10] ),
    .C(\top.compVal[9] ),
    .D(\top.compVal[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03396_));
 sky130_fd_sc_hd__or4_1 _06599_ (.A(\top.compVal[15] ),
    .B(\top.compVal[14] ),
    .C(\top.compVal[13] ),
    .D(\top.compVal[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03397_));
 sky130_fd_sc_hd__or4_1 _06600_ (.A(\top.compVal[7] ),
    .B(\top.compVal[6] ),
    .C(\top.compVal[5] ),
    .D(\top.compVal[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03398_));
 sky130_fd_sc_hd__or4_1 _06601_ (.A(\top.compVal[3] ),
    .B(\top.compVal[2] ),
    .C(\top.compVal[1] ),
    .D(\top.compVal[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03399_));
 sky130_fd_sc_hd__or4_1 _06602_ (.A(_03396_),
    .B(_03397_),
    .C(_03398_),
    .D(_03399_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03400_));
 sky130_fd_sc_hd__or4_1 _06603_ (.A(\top.compVal[27] ),
    .B(\top.compVal[26] ),
    .C(\top.compVal[25] ),
    .D(\top.compVal[24] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03401_));
 sky130_fd_sc_hd__or4_1 _06604_ (.A(\top.compVal[31] ),
    .B(\top.compVal[30] ),
    .C(\top.compVal[29] ),
    .D(\top.compVal[28] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03402_));
 sky130_fd_sc_hd__or4_1 _06605_ (.A(\top.compVal[23] ),
    .B(\top.compVal[22] ),
    .C(\top.compVal[21] ),
    .D(\top.compVal[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03403_));
 sky130_fd_sc_hd__or4_1 _06606_ (.A(\top.compVal[19] ),
    .B(\top.compVal[18] ),
    .C(\top.compVal[17] ),
    .D(\top.compVal[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03404_));
 sky130_fd_sc_hd__or3_1 _06607_ (.A(_03401_),
    .B(_03402_),
    .C(_03404_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03405_));
 sky130_fd_sc_hd__or4_1 _06608_ (.A(\top.compVal[43] ),
    .B(\top.compVal[42] ),
    .C(\top.compVal[41] ),
    .D(\top.compVal[40] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03406_));
 sky130_fd_sc_hd__or4_1 _06609_ (.A(\top.compVal[39] ),
    .B(\top.compVal[38] ),
    .C(\top.compVal[37] ),
    .D(\top.compVal[36] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03407_));
 sky130_fd_sc_hd__or4_1 _06610_ (.A(\top.compVal[35] ),
    .B(\top.compVal[34] ),
    .C(\top.compVal[33] ),
    .D(\top.compVal[32] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03408_));
 sky130_fd_sc_hd__or4_1 _06611_ (.A(\top.compVal[45] ),
    .B(\top.compVal[44] ),
    .C(_03406_),
    .D(_03408_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03409_));
 sky130_fd_sc_hd__or3_1 _06612_ (.A(_03400_),
    .B(_03407_),
    .C(_03409_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03410_));
 sky130_fd_sc_hd__or3_2 _06613_ (.A(_03403_),
    .B(_03405_),
    .C(_03410_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03411_));
 sky130_fd_sc_hd__and4b_2 _06614_ (.A_N(\top.controller.fin_FLV ),
    .B(_02500_),
    .C(net456),
    .D(_03411_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03412_));
 sky130_fd_sc_hd__and2_1 _06615_ (.A(_02429_),
    .B(\top.findLeastValue.val1[23] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03413_));
 sky130_fd_sc_hd__a22o_1 _06616_ (.A1(\top.compVal[21] ),
    .A2(_02492_),
    .B1(_02493_),
    .B2(\top.compVal[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03414_));
 sky130_fd_sc_hd__and2b_1 _06617_ (.A_N(\top.findLeastValue.val1[18] ),
    .B(\top.compVal[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03415_));
 sky130_fd_sc_hd__and2b_1 _06618_ (.A_N(\top.compVal[18] ),
    .B(\top.findLeastValue.val1[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03416_));
 sky130_fd_sc_hd__and2b_1 _06619_ (.A_N(\top.findLeastValue.val1[19] ),
    .B(\top.compVal[19] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03417_));
 sky130_fd_sc_hd__nand2b_1 _06620_ (.A_N(\top.compVal[19] ),
    .B(\top.findLeastValue.val1[19] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03418_));
 sky130_fd_sc_hd__or4b_1 _06621_ (.A(_03415_),
    .B(_03416_),
    .C(_03417_),
    .D_N(_03418_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03419_));
 sky130_fd_sc_hd__o22ai_1 _06622_ (.A1(_02432_),
    .A2(\top.findLeastValue.val1[17] ),
    .B1(\top.findLeastValue.val1[16] ),
    .B2(_02433_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03420_));
 sky130_fd_sc_hd__a21oi_1 _06623_ (.A1(_02432_),
    .A2(\top.findLeastValue.val1[17] ),
    .B1(_03419_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03421_));
 sky130_fd_sc_hd__a22o_1 _06624_ (.A1(_03415_),
    .A2(_03418_),
    .B1(_03420_),
    .B2(_03421_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03422_));
 sky130_fd_sc_hd__o22a_1 _06625_ (.A1(\top.compVal[20] ),
    .A2(_02493_),
    .B1(_03417_),
    .B2(_03422_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03423_));
 sky130_fd_sc_hd__o2bb2a_1 _06626_ (.A1_N(_02430_),
    .A2_N(\top.findLeastValue.val1[22] ),
    .B1(_02492_),
    .B2(\top.compVal[21] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03424_));
 sky130_fd_sc_hd__o21ai_1 _06627_ (.A1(_03414_),
    .A2(_03423_),
    .B1(_03424_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03425_));
 sky130_fd_sc_hd__o221ai_1 _06628_ (.A1(_02429_),
    .A2(\top.findLeastValue.val1[23] ),
    .B1(\top.findLeastValue.val1[22] ),
    .B2(_02430_),
    .C1(_03424_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03426_));
 sky130_fd_sc_hd__o221a_1 _06629_ (.A1(_02429_),
    .A2(\top.findLeastValue.val1[23] ),
    .B1(\top.findLeastValue.val1[22] ),
    .B2(_02430_),
    .C1(_03425_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03427_));
 sky130_fd_sc_hd__a2bb2o_1 _06630_ (.A1_N(_02434_),
    .A2_N(\top.findLeastValue.val1[15] ),
    .B1(_02494_),
    .B2(\top.compVal[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03428_));
 sky130_fd_sc_hd__and2b_1 _06631_ (.A_N(\top.findLeastValue.val1[12] ),
    .B(\top.compVal[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03429_));
 sky130_fd_sc_hd__and2_1 _06632_ (.A(_02439_),
    .B(\top.findLeastValue.val1[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03430_));
 sky130_fd_sc_hd__o22a_1 _06633_ (.A1(_02441_),
    .A2(\top.findLeastValue.val1[5] ),
    .B1(\top.findLeastValue.val1[4] ),
    .B2(_02442_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03431_));
 sky130_fd_sc_hd__o22a_1 _06634_ (.A1(_02443_),
    .A2(\top.findLeastValue.val1[3] ),
    .B1(\top.findLeastValue.val1[2] ),
    .B2(_02444_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03432_));
 sky130_fd_sc_hd__o211a_1 _06635_ (.A1(_02445_),
    .A2(\top.findLeastValue.val1[1] ),
    .B1(\top.findLeastValue.val1[0] ),
    .C1(_02446_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03433_));
 sky130_fd_sc_hd__a22o_1 _06636_ (.A1(_02444_),
    .A2(\top.findLeastValue.val1[2] ),
    .B1(\top.findLeastValue.val1[1] ),
    .B2(_02445_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03434_));
 sky130_fd_sc_hd__o21a_1 _06637_ (.A1(_03433_),
    .A2(_03434_),
    .B1(_03432_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03435_));
 sky130_fd_sc_hd__and2_1 _06638_ (.A(_02442_),
    .B(\top.findLeastValue.val1[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03436_));
 sky130_fd_sc_hd__nor2_1 _06639_ (.A(\top.compVal[5] ),
    .B(_02498_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03437_));
 sky130_fd_sc_hd__o22ai_1 _06640_ (.A1(_02439_),
    .A2(\top.findLeastValue.val1[7] ),
    .B1(\top.findLeastValue.val1[6] ),
    .B2(_02440_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03438_));
 sky130_fd_sc_hd__nand2b_1 _06641_ (.A_N(_03430_),
    .B(_03438_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03439_));
 sky130_fd_sc_hd__a211o_1 _06642_ (.A1(_02440_),
    .A2(\top.findLeastValue.val1[6] ),
    .B1(_03430_),
    .C1(_03438_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03440_));
 sky130_fd_sc_hd__or3_1 _06643_ (.A(_03431_),
    .B(_03437_),
    .C(_03440_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03441_));
 sky130_fd_sc_hd__or3b_1 _06644_ (.A(_03436_),
    .B(_03437_),
    .C_N(_03431_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03442_));
 sky130_fd_sc_hd__a2111o_1 _06645_ (.A1(_02443_),
    .A2(\top.findLeastValue.val1[3] ),
    .B1(_03435_),
    .C1(_03440_),
    .D1(_03442_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03443_));
 sky130_fd_sc_hd__a32o_1 _06646_ (.A1(_03439_),
    .A2(_03441_),
    .A3(_03443_),
    .B1(\top.findLeastValue.val1[8] ),
    .B2(_02438_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03444_));
 sky130_fd_sc_hd__o221a_1 _06647_ (.A1(_02437_),
    .A2(\top.findLeastValue.val1[9] ),
    .B1(\top.findLeastValue.val1[8] ),
    .B2(_02438_),
    .C1(_03444_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03445_));
 sky130_fd_sc_hd__o22a_1 _06648_ (.A1(_02435_),
    .A2(\top.findLeastValue.val1[11] ),
    .B1(\top.findLeastValue.val1[10] ),
    .B2(_02436_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03446_));
 sky130_fd_sc_hd__and2_1 _06649_ (.A(_02435_),
    .B(\top.findLeastValue.val1[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03447_));
 sky130_fd_sc_hd__a22o_1 _06650_ (.A1(_02436_),
    .A2(\top.findLeastValue.val1[10] ),
    .B1(\top.findLeastValue.val1[9] ),
    .B2(_02437_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03448_));
 sky130_fd_sc_hd__or3b_1 _06651_ (.A(_03447_),
    .B(_03448_),
    .C_N(_03446_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03449_));
 sky130_fd_sc_hd__o22ai_1 _06652_ (.A1(_03446_),
    .A2(_03447_),
    .B1(_03449_),
    .B2(_03445_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03450_));
 sky130_fd_sc_hd__nand2b_1 _06653_ (.A_N(\top.compVal[12] ),
    .B(\top.findLeastValue.val1[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03451_));
 sky130_fd_sc_hd__a221o_1 _06654_ (.A1(\top.compVal[13] ),
    .A2(_02495_),
    .B1(_03450_),
    .B2(_03451_),
    .C1(_03429_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03452_));
 sky130_fd_sc_hd__o22a_1 _06655_ (.A1(\top.compVal[14] ),
    .A2(_02494_),
    .B1(_02495_),
    .B2(\top.compVal[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03453_));
 sky130_fd_sc_hd__a21oi_1 _06656_ (.A1(_03452_),
    .A2(_03453_),
    .B1(_03428_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03454_));
 sky130_fd_sc_hd__a211o_1 _06657_ (.A1(_02434_),
    .A2(\top.findLeastValue.val1[15] ),
    .B1(_03413_),
    .C1(_03420_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03455_));
 sky130_fd_sc_hd__a221o_1 _06658_ (.A1(_02432_),
    .A2(\top.findLeastValue.val1[17] ),
    .B1(\top.findLeastValue.val1[16] ),
    .B2(_02433_),
    .C1(_03455_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03456_));
 sky130_fd_sc_hd__a2111o_1 _06659_ (.A1(_02431_),
    .A2(\top.findLeastValue.val1[20] ),
    .B1(_03414_),
    .C1(_03419_),
    .D1(_03456_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03457_));
 sky130_fd_sc_hd__o32a_1 _06660_ (.A1(_03426_),
    .A2(_03454_),
    .A3(_03457_),
    .B1(_03427_),
    .B2(_03413_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03458_));
 sky130_fd_sc_hd__a22o_1 _06661_ (.A1(_02423_),
    .A2(\top.findLeastValue.val1[29] ),
    .B1(\top.findLeastValue.val1[28] ),
    .B2(_02424_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03459_));
 sky130_fd_sc_hd__a22o_1 _06662_ (.A1(\top.compVal[27] ),
    .A2(_02490_),
    .B1(\top.findLeastValue.val1[26] ),
    .B2(_02426_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03460_));
 sky130_fd_sc_hd__o22a_1 _06663_ (.A1(_02427_),
    .A2(\top.findLeastValue.val1[25] ),
    .B1(\top.findLeastValue.val1[24] ),
    .B2(_02428_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03461_));
 sky130_fd_sc_hd__o22ai_2 _06664_ (.A1(_02422_),
    .A2(\top.findLeastValue.val1[30] ),
    .B1(\top.findLeastValue.val1[29] ),
    .B2(_02423_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03462_));
 sky130_fd_sc_hd__nor2_1 _06665_ (.A(\top.compVal[27] ),
    .B(_02490_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03463_));
 sky130_fd_sc_hd__a22o_1 _06666_ (.A1(_02421_),
    .A2(\top.findLeastValue.val1[31] ),
    .B1(\top.findLeastValue.val1[30] ),
    .B2(_02422_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03464_));
 sky130_fd_sc_hd__or2_1 _06667_ (.A(_02421_),
    .B(\top.findLeastValue.val1[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03465_));
 sky130_fd_sc_hd__and2_1 _06668_ (.A(_02427_),
    .B(\top.findLeastValue.val1[25] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03466_));
 sky130_fd_sc_hd__a2bb2o_1 _06669_ (.A1_N(_02424_),
    .A2_N(\top.findLeastValue.val1[28] ),
    .B1(\top.findLeastValue.val1[24] ),
    .B2(_02428_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03467_));
 sky130_fd_sc_hd__or4_1 _06670_ (.A(_03459_),
    .B(_03460_),
    .C(_03462_),
    .D(_03464_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03468_));
 sky130_fd_sc_hd__a2111oi_1 _06671_ (.A1(\top.compVal[26] ),
    .A2(_02491_),
    .B1(_03466_),
    .C1(_03467_),
    .D1(_03468_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03469_));
 sky130_fd_sc_hd__nand2_1 _06672_ (.A(_03461_),
    .B(_03469_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03470_));
 sky130_fd_sc_hd__o32a_1 _06673_ (.A1(_03460_),
    .A2(_03461_),
    .A3(_03466_),
    .B1(\top.findLeastValue.val1[26] ),
    .B2(_02426_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03471_));
 sky130_fd_sc_hd__or2_1 _06674_ (.A(_03463_),
    .B(_03471_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03472_));
 sky130_fd_sc_hd__o221a_1 _06675_ (.A1(_02424_),
    .A2(\top.findLeastValue.val1[28] ),
    .B1(\top.findLeastValue.val1[27] ),
    .B2(_02425_),
    .C1(_03472_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03473_));
 sky130_fd_sc_hd__nor2_1 _06676_ (.A(_03459_),
    .B(_03473_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03474_));
 sky130_fd_sc_hd__o21bai_2 _06677_ (.A1(_03462_),
    .A2(_03474_),
    .B1_N(_03464_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03475_));
 sky130_fd_sc_hd__o311ai_4 _06678_ (.A1(_03458_),
    .A2(_03463_),
    .A3(_03470_),
    .B1(_03475_),
    .C1(_03465_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03476_));
 sky130_fd_sc_hd__a22o_1 _06679_ (.A1(\top.compVal[41] ),
    .A2(_02482_),
    .B1(_02483_),
    .B2(\top.compVal[40] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03477_));
 sky130_fd_sc_hd__a22o_1 _06680_ (.A1(\top.compVal[33] ),
    .A2(_02488_),
    .B1(_02489_),
    .B2(\top.compVal[32] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03478_));
 sky130_fd_sc_hd__a22o_1 _06681_ (.A1(_02410_),
    .A2(\top.findLeastValue.val1[37] ),
    .B1(\top.findLeastValue.val1[36] ),
    .B2(_02411_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03479_));
 sky130_fd_sc_hd__o22a_1 _06682_ (.A1(\top.compVal[40] ),
    .A2(_02483_),
    .B1(_02484_),
    .B2(\top.compVal[39] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03480_));
 sky130_fd_sc_hd__and2_1 _06683_ (.A(\top.compVal[39] ),
    .B(_02484_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03481_));
 sky130_fd_sc_hd__a221o_1 _06684_ (.A1(\top.compVal[38] ),
    .A2(_02485_),
    .B1(_02486_),
    .B2(\top.compVal[37] ),
    .C1(_03481_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03482_));
 sky130_fd_sc_hd__nand2_1 _06685_ (.A(_02414_),
    .B(\top.findLeastValue.val1[33] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03483_));
 sky130_fd_sc_hd__a21o_1 _06686_ (.A1(_02406_),
    .A2(\top.findLeastValue.val1[45] ),
    .B1(\top.findLeastValue.val1[46] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03484_));
 sky130_fd_sc_hd__o22a_1 _06687_ (.A1(_02406_),
    .A2(\top.findLeastValue.val1[45] ),
    .B1(\top.findLeastValue.val1[44] ),
    .B2(_02407_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03485_));
 sky130_fd_sc_hd__a21oi_1 _06688_ (.A1(_02408_),
    .A2(\top.findLeastValue.val1[43] ),
    .B1(_03484_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03486_));
 sky130_fd_sc_hd__o211a_1 _06689_ (.A1(\top.compVal[44] ),
    .A2(_02480_),
    .B1(_03485_),
    .C1(_03486_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03487_));
 sky130_fd_sc_hd__o221a_1 _06690_ (.A1(\top.compVal[42] ),
    .A2(_02481_),
    .B1(_02482_),
    .B2(\top.compVal[41] ),
    .C1(_03487_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03488_));
 sky130_fd_sc_hd__inv_2 _06691_ (.A(_03488_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03489_));
 sky130_fd_sc_hd__a2bb2o_1 _06692_ (.A1_N(_02408_),
    .A2_N(\top.findLeastValue.val1[43] ),
    .B1(_02481_),
    .B2(\top.compVal[42] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03490_));
 sky130_fd_sc_hd__o22a_1 _06693_ (.A1(_02411_),
    .A2(\top.findLeastValue.val1[36] ),
    .B1(\top.findLeastValue.val1[35] ),
    .B2(_02412_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03491_));
 sky130_fd_sc_hd__a22o_1 _06694_ (.A1(_02412_),
    .A2(\top.findLeastValue.val1[35] ),
    .B1(\top.findLeastValue.val1[34] ),
    .B2(_02413_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03492_));
 sky130_fd_sc_hd__nand2b_1 _06695_ (.A_N(_03479_),
    .B(_03491_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03493_));
 sky130_fd_sc_hd__a221o_1 _06696_ (.A1(_02409_),
    .A2(\top.findLeastValue.val1[38] ),
    .B1(\top.findLeastValue.val1[33] ),
    .B2(_02414_),
    .C1(_03492_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03494_));
 sky130_fd_sc_hd__or4_1 _06697_ (.A(_03477_),
    .B(_03482_),
    .C(_03493_),
    .D(_03494_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03495_));
 sky130_fd_sc_hd__o221a_1 _06698_ (.A1(_02413_),
    .A2(\top.findLeastValue.val1[34] ),
    .B1(_02489_),
    .B2(\top.compVal[32] ),
    .C1(_03480_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03496_));
 sky130_fd_sc_hd__or4b_1 _06699_ (.A(_03478_),
    .B(_03489_),
    .C(_03490_),
    .D_N(_03496_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03497_));
 sky130_fd_sc_hd__nor2_1 _06700_ (.A(_03495_),
    .B(_03497_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03498_));
 sky130_fd_sc_hd__o2bb2a_1 _06701_ (.A1_N(_03478_),
    .A2_N(_03483_),
    .B1(_02413_),
    .B2(\top.findLeastValue.val1[34] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03499_));
 sky130_fd_sc_hd__o21a_1 _06702_ (.A1(_03492_),
    .A2(_03499_),
    .B1(_03491_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03500_));
 sky130_fd_sc_hd__o21bai_1 _06703_ (.A1(_03479_),
    .A2(_03500_),
    .B1_N(_03482_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03501_));
 sky130_fd_sc_hd__o311a_1 _06704_ (.A1(\top.compVal[38] ),
    .A2(_02485_),
    .A3(_03481_),
    .B1(_03501_),
    .C1(_03480_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03502_));
 sky130_fd_sc_hd__o21ai_1 _06705_ (.A1(_03477_),
    .A2(_03502_),
    .B1(_03488_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03503_));
 sky130_fd_sc_hd__o2bb2a_1 _06706_ (.A1_N(_03490_),
    .A2_N(_03487_),
    .B1(_03485_),
    .B2(_03484_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03504_));
 sky130_fd_sc_hd__nand2_1 _06707_ (.A(_03503_),
    .B(_03504_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03505_));
 sky130_fd_sc_hd__a21oi_1 _06708_ (.A1(_03476_),
    .A2(_03498_),
    .B1(_03505_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03506_));
 sky130_fd_sc_hd__a21oi_1 _06709_ (.A1(_03412_),
    .A2(net149),
    .B1(net288),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03507_));
 sky130_fd_sc_hd__a21o_1 _06710_ (.A1(_03412_),
    .A2(net149),
    .B1(net288),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03508_));
 sky130_fd_sc_hd__a2bb2o_1 _06711_ (.A1_N(_02406_),
    .A2_N(\top.findLeastValue.val2[45] ),
    .B1(_02455_),
    .B2(\top.compVal[44] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03509_));
 sky130_fd_sc_hd__a22o_1 _06712_ (.A1(\top.compVal[41] ),
    .A2(_02457_),
    .B1(_02458_),
    .B2(\top.compVal[40] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03510_));
 sky130_fd_sc_hd__o22a_1 _06713_ (.A1(\top.compVal[42] ),
    .A2(_02456_),
    .B1(_02457_),
    .B2(\top.compVal[41] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03511_));
 sky130_fd_sc_hd__nand2_1 _06714_ (.A(_03510_),
    .B(_03511_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03512_));
 sky130_fd_sc_hd__o2bb2a_1 _06715_ (.A1_N(_02456_),
    .A2_N(\top.compVal[42] ),
    .B1(_02408_),
    .B2(\top.findLeastValue.val2[43] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03513_));
 sky130_fd_sc_hd__a22o_1 _06716_ (.A1(_02407_),
    .A2(\top.findLeastValue.val2[44] ),
    .B1(\top.findLeastValue.val2[43] ),
    .B2(_02408_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03514_));
 sky130_fd_sc_hd__a21oi_1 _06717_ (.A1(_03512_),
    .A2(_03513_),
    .B1(_03514_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03515_));
 sky130_fd_sc_hd__a2bb2o_1 _06718_ (.A1_N(_03509_),
    .A2_N(_03515_),
    .B1(_02406_),
    .B2(\top.findLeastValue.val2[45] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03516_));
 sky130_fd_sc_hd__nand2_1 _06719_ (.A(_02409_),
    .B(\top.findLeastValue.val2[38] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03517_));
 sky130_fd_sc_hd__nand2_1 _06720_ (.A(_02414_),
    .B(\top.findLeastValue.val2[33] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03518_));
 sky130_fd_sc_hd__and3b_1 _06721_ (.A_N(\top.findLeastValue.val2[32] ),
    .B(_03518_),
    .C(\top.compVal[32] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03519_));
 sky130_fd_sc_hd__a221o_1 _06722_ (.A1(\top.compVal[34] ),
    .A2(_02463_),
    .B1(_02464_),
    .B2(\top.compVal[33] ),
    .C1(_03519_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03520_));
 sky130_fd_sc_hd__o22a_1 _06723_ (.A1(\top.compVal[37] ),
    .A2(_02460_),
    .B1(_02461_),
    .B2(\top.compVal[36] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03521_));
 sky130_fd_sc_hd__o22a_1 _06724_ (.A1(\top.compVal[35] ),
    .A2(_02462_),
    .B1(_02463_),
    .B2(\top.compVal[34] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03522_));
 sky130_fd_sc_hd__and3_1 _06725_ (.A(_03520_),
    .B(_03521_),
    .C(_03522_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03523_));
 sky130_fd_sc_hd__a22o_1 _06726_ (.A1(\top.compVal[36] ),
    .A2(_02461_),
    .B1(_02462_),
    .B2(\top.compVal[35] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03524_));
 sky130_fd_sc_hd__a22o_1 _06727_ (.A1(\top.compVal[37] ),
    .A2(_02460_),
    .B1(_03521_),
    .B2(_03524_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03525_));
 sky130_fd_sc_hd__o21a_1 _06728_ (.A1(_03523_),
    .A2(_03525_),
    .B1(_03517_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03526_));
 sky130_fd_sc_hd__a2bb2o_1 _06729_ (.A1_N(\top.findLeastValue.val2[38] ),
    .A2_N(_02409_),
    .B1(\top.compVal[39] ),
    .B2(_02459_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03527_));
 sky130_fd_sc_hd__nand2_1 _06730_ (.A(_02435_),
    .B(\top.findLeastValue.val2[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03528_));
 sky130_fd_sc_hd__a2bb2o_1 _06731_ (.A1_N(_02435_),
    .A2_N(\top.findLeastValue.val2[11] ),
    .B1(_02474_),
    .B2(\top.compVal[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03529_));
 sky130_fd_sc_hd__a21oi_1 _06732_ (.A1(_02436_),
    .A2(\top.findLeastValue.val2[10] ),
    .B1(_03529_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03530_));
 sky130_fd_sc_hd__o211a_1 _06733_ (.A1(\top.compVal[9] ),
    .A2(_02475_),
    .B1(_03528_),
    .C1(_03530_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03531_));
 sky130_fd_sc_hd__a22o_1 _06734_ (.A1(\top.compVal[9] ),
    .A2(_02475_),
    .B1(_02476_),
    .B2(\top.compVal[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03532_));
 sky130_fd_sc_hd__and2b_1 _06735_ (.A_N(\top.findLeastValue.val2[1] ),
    .B(\top.compVal[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03533_));
 sky130_fd_sc_hd__nand2b_1 _06736_ (.A_N(\top.compVal[2] ),
    .B(\top.findLeastValue.val2[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03534_));
 sky130_fd_sc_hd__nand2b_1 _06737_ (.A_N(\top.compVal[1] ),
    .B(\top.findLeastValue.val2[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03535_));
 sky130_fd_sc_hd__o311a_1 _06738_ (.A1(\top.compVal[0] ),
    .A2(_02479_),
    .A3(_03533_),
    .B1(_03534_),
    .C1(_03535_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03536_));
 sky130_fd_sc_hd__a2bb2o_1 _06739_ (.A1_N(\top.findLeastValue.val2[2] ),
    .A2_N(_02444_),
    .B1(\top.compVal[3] ),
    .B2(_02478_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03537_));
 sky130_fd_sc_hd__nand2_1 _06740_ (.A(_02442_),
    .B(\top.findLeastValue.val2[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03538_));
 sky130_fd_sc_hd__o221a_1 _06741_ (.A1(\top.compVal[3] ),
    .A2(_02478_),
    .B1(_03536_),
    .B2(_03537_),
    .C1(_03538_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03539_));
 sky130_fd_sc_hd__a2bb2o_1 _06742_ (.A1_N(\top.findLeastValue.val2[4] ),
    .A2_N(_02442_),
    .B1(\top.compVal[5] ),
    .B2(_02477_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03540_));
 sky130_fd_sc_hd__a22o_1 _06743_ (.A1(_02440_),
    .A2(\top.findLeastValue.val2[6] ),
    .B1(\top.findLeastValue.val2[5] ),
    .B2(_02441_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03541_));
 sky130_fd_sc_hd__o21bai_1 _06744_ (.A1(_03539_),
    .A2(_03540_),
    .B1_N(_03541_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03542_));
 sky130_fd_sc_hd__o22a_1 _06745_ (.A1(_02439_),
    .A2(\top.findLeastValue.val2[7] ),
    .B1(\top.findLeastValue.val2[6] ),
    .B2(_02440_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03543_));
 sky130_fd_sc_hd__a22o_1 _06746_ (.A1(_03528_),
    .A2(_03529_),
    .B1(_03531_),
    .B2(_03532_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03544_));
 sky130_fd_sc_hd__a221o_1 _06747_ (.A1(_02438_),
    .A2(\top.findLeastValue.val2[8] ),
    .B1(\top.findLeastValue.val2[7] ),
    .B2(_02439_),
    .C1(_03532_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03545_));
 sky130_fd_sc_hd__a21oi_1 _06748_ (.A1(_03542_),
    .A2(_03543_),
    .B1(_03545_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03546_));
 sky130_fd_sc_hd__a21o_1 _06749_ (.A1(_03531_),
    .A2(_03546_),
    .B1(_03544_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03547_));
 sky130_fd_sc_hd__nor2_1 _06750_ (.A(_02434_),
    .B(\top.findLeastValue.val2[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03548_));
 sky130_fd_sc_hd__a2bb2o_1 _06751_ (.A1_N(_02472_),
    .A2_N(\top.compVal[14] ),
    .B1(_02434_),
    .B2(\top.findLeastValue.val2[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03549_));
 sky130_fd_sc_hd__a211o_1 _06752_ (.A1(\top.compVal[14] ),
    .A2(_02472_),
    .B1(_03548_),
    .C1(_03549_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03550_));
 sky130_fd_sc_hd__and2_1 _06753_ (.A(\top.compVal[13] ),
    .B(_02473_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03551_));
 sky130_fd_sc_hd__or2_1 _06754_ (.A(\top.compVal[13] ),
    .B(_02473_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03552_));
 sky130_fd_sc_hd__xor2_1 _06755_ (.A(\top.compVal[12] ),
    .B(\top.findLeastValue.val2[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03553_));
 sky130_fd_sc_hd__nor3_1 _06756_ (.A(_03550_),
    .B(_03551_),
    .C(_03553_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03554_));
 sky130_fd_sc_hd__and3b_1 _06757_ (.A_N(\top.findLeastValue.val2[12] ),
    .B(_03552_),
    .C(\top.compVal[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03555_));
 sky130_fd_sc_hd__o21ba_1 _06758_ (.A1(_03551_),
    .A2(_03555_),
    .B1_N(_03550_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03556_));
 sky130_fd_sc_hd__a21oi_1 _06759_ (.A1(_02434_),
    .A2(\top.findLeastValue.val2[15] ),
    .B1(\top.findLeastValue.val2[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03557_));
 sky130_fd_sc_hd__a211o_1 _06760_ (.A1(\top.compVal[14] ),
    .A2(_03557_),
    .B1(_03556_),
    .C1(_03548_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03558_));
 sky130_fd_sc_hd__a31o_1 _06761_ (.A1(_03547_),
    .A2(_03552_),
    .A3(_03554_),
    .B1(_03558_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03559_));
 sky130_fd_sc_hd__and2_1 _06762_ (.A(\top.compVal[19] ),
    .B(_02469_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03560_));
 sky130_fd_sc_hd__nand2_1 _06763_ (.A(_02432_),
    .B(\top.findLeastValue.val2[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03561_));
 sky130_fd_sc_hd__a2bb2o_1 _06764_ (.A1_N(\top.findLeastValue.val2[17] ),
    .A2_N(_02432_),
    .B1(\top.compVal[18] ),
    .B2(_02470_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03562_));
 sky130_fd_sc_hd__a221o_1 _06765_ (.A1(_02432_),
    .A2(\top.findLeastValue.val2[17] ),
    .B1(_02471_),
    .B2(\top.compVal[16] ),
    .C1(_03562_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03563_));
 sky130_fd_sc_hd__nand2b_1 _06766_ (.A_N(\top.findLeastValue.val2[21] ),
    .B(\top.compVal[21] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03564_));
 sky130_fd_sc_hd__a22o_1 _06767_ (.A1(\top.compVal[29] ),
    .A2(_02465_),
    .B1(_02466_),
    .B2(\top.compVal[28] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03565_));
 sky130_fd_sc_hd__inv_2 _06768_ (.A(_03565_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03566_));
 sky130_fd_sc_hd__o22a_1 _06769_ (.A1(_02427_),
    .A2(\top.findLeastValue.val2[25] ),
    .B1(\top.findLeastValue.val2[24] ),
    .B2(_02428_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03567_));
 sky130_fd_sc_hd__o22a_1 _06770_ (.A1(_02425_),
    .A2(\top.findLeastValue.val2[27] ),
    .B1(\top.findLeastValue.val2[26] ),
    .B2(_02426_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03568_));
 sky130_fd_sc_hd__nand2_1 _06771_ (.A(_02425_),
    .B(\top.findLeastValue.val2[27] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03569_));
 sky130_fd_sc_hd__nand2_1 _06772_ (.A(_02427_),
    .B(\top.findLeastValue.val2[25] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03570_));
 sky130_fd_sc_hd__o211a_1 _06773_ (.A1(\top.compVal[26] ),
    .A2(_02467_),
    .B1(_03568_),
    .C1(_03569_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03571_));
 sky130_fd_sc_hd__o22a_1 _06774_ (.A1(_02421_),
    .A2(\top.findLeastValue.val2[31] ),
    .B1(\top.findLeastValue.val2[30] ),
    .B2(_02422_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03572_));
 sky130_fd_sc_hd__a22oi_1 _06775_ (.A1(_02421_),
    .A2(\top.findLeastValue.val2[31] ),
    .B1(\top.findLeastValue.val2[30] ),
    .B2(_02422_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03573_));
 sky130_fd_sc_hd__o211a_1 _06776_ (.A1(\top.compVal[29] ),
    .A2(_02465_),
    .B1(_03572_),
    .C1(_03573_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03574_));
 sky130_fd_sc_hd__xnor2_1 _06777_ (.A(\top.compVal[22] ),
    .B(\top.findLeastValue.val2[22] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03575_));
 sky130_fd_sc_hd__nand2b_1 _06778_ (.A_N(\top.compVal[23] ),
    .B(\top.findLeastValue.val2[23] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03576_));
 sky130_fd_sc_hd__nand2b_1 _06779_ (.A_N(\top.findLeastValue.val2[23] ),
    .B(\top.compVal[23] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03577_));
 sky130_fd_sc_hd__nand2b_1 _06780_ (.A_N(\top.compVal[21] ),
    .B(\top.findLeastValue.val2[21] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03578_));
 sky130_fd_sc_hd__o2111a_1 _06781_ (.A1(\top.compVal[24] ),
    .A2(_02468_),
    .B1(_03567_),
    .C1(_03570_),
    .D1(_03571_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03579_));
 sky130_fd_sc_hd__and3_1 _06782_ (.A(_03575_),
    .B(_03576_),
    .C(_03577_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03580_));
 sky130_fd_sc_hd__xnor2_1 _06783_ (.A(\top.compVal[20] ),
    .B(\top.findLeastValue.val2[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03581_));
 sky130_fd_sc_hd__o211a_1 _06784_ (.A1(\top.compVal[28] ),
    .A2(_02466_),
    .B1(_03566_),
    .C1(_03574_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03582_));
 sky130_fd_sc_hd__and4_1 _06785_ (.A(_03564_),
    .B(_03578_),
    .C(_03580_),
    .D(_03581_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03583_));
 sky130_fd_sc_hd__and3_1 _06786_ (.A(_03579_),
    .B(_03582_),
    .C(_03583_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03584_));
 sky130_fd_sc_hd__o221ai_1 _06787_ (.A1(\top.compVal[19] ),
    .A2(_02469_),
    .B1(_02470_),
    .B2(\top.compVal[18] ),
    .C1(_03584_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03585_));
 sky130_fd_sc_hd__a2111oi_1 _06788_ (.A1(_02433_),
    .A2(\top.findLeastValue.val2[16] ),
    .B1(_03560_),
    .C1(_03563_),
    .D1(_03585_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03586_));
 sky130_fd_sc_hd__and2b_1 _06789_ (.A_N(_03568_),
    .B(_03569_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03587_));
 sky130_fd_sc_hd__or3b_1 _06790_ (.A(_02431_),
    .B(\top.findLeastValue.val2[20] ),
    .C_N(_03578_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03588_));
 sky130_fd_sc_hd__a21bo_1 _06791_ (.A1(_03564_),
    .A2(_03588_),
    .B1_N(_03580_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03589_));
 sky130_fd_sc_hd__or3b_1 _06792_ (.A(_02430_),
    .B(\top.findLeastValue.val2[22] ),
    .C_N(_03576_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03590_));
 sky130_fd_sc_hd__a32o_1 _06793_ (.A1(_03577_),
    .A2(_03589_),
    .A3(_03590_),
    .B1(\top.findLeastValue.val2[24] ),
    .B2(_02428_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03591_));
 sky130_fd_sc_hd__nand2_1 _06794_ (.A(_03567_),
    .B(_03591_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03592_));
 sky130_fd_sc_hd__a31o_1 _06795_ (.A1(_03570_),
    .A2(_03571_),
    .A3(_03592_),
    .B1(_03587_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03593_));
 sky130_fd_sc_hd__a31o_1 _06796_ (.A1(\top.compVal[16] ),
    .A2(_02471_),
    .A3(_03561_),
    .B1(_03562_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03594_));
 sky130_fd_sc_hd__a21oi_1 _06797_ (.A1(_02421_),
    .A2(\top.findLeastValue.val2[31] ),
    .B1(_03572_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03595_));
 sky130_fd_sc_hd__o221a_1 _06798_ (.A1(\top.compVal[19] ),
    .A2(_02469_),
    .B1(_02470_),
    .B2(\top.compVal[18] ),
    .C1(_03594_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03596_));
 sky130_fd_sc_hd__o21a_1 _06799_ (.A1(_03560_),
    .A2(_03596_),
    .B1(_03584_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03597_));
 sky130_fd_sc_hd__a221o_1 _06800_ (.A1(_03565_),
    .A2(_03574_),
    .B1(_03582_),
    .B2(_03593_),
    .C1(_03597_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03598_));
 sky130_fd_sc_hd__a211o_1 _06801_ (.A1(_03559_),
    .A2(_03586_),
    .B1(_03595_),
    .C1(_03598_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03599_));
 sky130_fd_sc_hd__o221a_1 _06802_ (.A1(_02411_),
    .A2(\top.findLeastValue.val2[36] ),
    .B1(\top.findLeastValue.val2[35] ),
    .B2(_02412_),
    .C1(_03521_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03600_));
 sky130_fd_sc_hd__o221a_1 _06803_ (.A1(_02413_),
    .A2(\top.findLeastValue.val2[34] ),
    .B1(\top.findLeastValue.val2[33] ),
    .B2(_02414_),
    .C1(_03522_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03601_));
 sky130_fd_sc_hd__o2bb2a_1 _06804_ (.A1_N(_02415_),
    .A2_N(\top.findLeastValue.val2[32] ),
    .B1(\top.findLeastValue.val2[37] ),
    .B2(_02410_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03602_));
 sky130_fd_sc_hd__o2111a_1 _06805_ (.A1(_02415_),
    .A2(\top.findLeastValue.val2[32] ),
    .B1(_03517_),
    .C1(_03518_),
    .D1(_03602_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03603_));
 sky130_fd_sc_hd__and4_1 _06806_ (.A(_03599_),
    .B(_03600_),
    .C(_03601_),
    .D(_03603_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03604_));
 sky130_fd_sc_hd__o32a_1 _06807_ (.A1(_03526_),
    .A2(_03527_),
    .A3(_03604_),
    .B1(_02459_),
    .B2(\top.compVal[39] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03605_));
 sky130_fd_sc_hd__o21bai_1 _06808_ (.A1(\top.compVal[40] ),
    .A2(_02458_),
    .B1_N(_03514_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03606_));
 sky130_fd_sc_hd__a2111oi_1 _06809_ (.A1(_02406_),
    .A2(\top.findLeastValue.val2[45] ),
    .B1(_03509_),
    .C1(_03606_),
    .D1(\top.findLeastValue.val2[46] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03607_));
 sky130_fd_sc_hd__and4b_1 _06810_ (.A_N(_03510_),
    .B(_03511_),
    .C(_03513_),
    .D(_03607_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03608_));
 sky130_fd_sc_hd__o2bb2a_2 _06811_ (.A1_N(_03608_),
    .A2_N(_03605_),
    .B1(_03516_),
    .B2(\top.findLeastValue.val2[46] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03609_));
 sky130_fd_sc_hd__and2_1 _06812_ (.A(_03412_),
    .B(_03609_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03610_));
 sky130_fd_sc_hd__a211o_1 _06813_ (.A1(_03412_),
    .A2(net149),
    .B1(_03610_),
    .C1(net288),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03611_));
 sky130_fd_sc_hd__and2_1 _06814_ (.A(net287),
    .B(net125),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03612_));
 sky130_fd_sc_hd__nand2_1 _06815_ (.A(_03394_),
    .B(net126),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03613_));
 sky130_fd_sc_hd__o22a_1 _06816_ (.A1(\top.findLeastValue.val2[46] ),
    .A2(net128),
    .B1(net119),
    .B2(\top.findLeastValue.val1[46] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02054_));
 sky130_fd_sc_hd__mux2_1 _06817_ (.A0(\top.compVal[45] ),
    .A1(\top.findLeastValue.val1[45] ),
    .S(net152),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03614_));
 sky130_fd_sc_hd__o22a_1 _06818_ (.A1(\top.findLeastValue.val2[45] ),
    .A2(net131),
    .B1(net119),
    .B2(_03614_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02053_));
 sky130_fd_sc_hd__mux2_1 _06819_ (.A0(\top.compVal[44] ),
    .A1(\top.findLeastValue.val1[44] ),
    .S(net153),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03615_));
 sky130_fd_sc_hd__o22a_1 _06820_ (.A1(\top.findLeastValue.val2[44] ),
    .A2(net129),
    .B1(net119),
    .B2(_03615_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02052_));
 sky130_fd_sc_hd__mux2_1 _06821_ (.A0(\top.compVal[43] ),
    .A1(\top.findLeastValue.val1[43] ),
    .S(net153),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03616_));
 sky130_fd_sc_hd__o22a_1 _06822_ (.A1(\top.findLeastValue.val2[43] ),
    .A2(net129),
    .B1(net119),
    .B2(_03616_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02051_));
 sky130_fd_sc_hd__mux2_1 _06823_ (.A0(\top.compVal[42] ),
    .A1(\top.findLeastValue.val1[42] ),
    .S(net153),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03617_));
 sky130_fd_sc_hd__o22a_1 _06824_ (.A1(\top.findLeastValue.val2[42] ),
    .A2(net129),
    .B1(net119),
    .B2(_03617_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02050_));
 sky130_fd_sc_hd__mux2_1 _06825_ (.A0(\top.compVal[41] ),
    .A1(\top.findLeastValue.val1[41] ),
    .S(net153),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03618_));
 sky130_fd_sc_hd__o22a_1 _06826_ (.A1(\top.findLeastValue.val2[41] ),
    .A2(net129),
    .B1(net119),
    .B2(_03618_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02049_));
 sky130_fd_sc_hd__mux2_1 _06827_ (.A0(\top.compVal[40] ),
    .A1(\top.findLeastValue.val1[40] ),
    .S(net153),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03619_));
 sky130_fd_sc_hd__o22a_1 _06828_ (.A1(\top.findLeastValue.val2[40] ),
    .A2(net129),
    .B1(net119),
    .B2(_03619_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02048_));
 sky130_fd_sc_hd__mux2_1 _06829_ (.A0(\top.compVal[39] ),
    .A1(\top.findLeastValue.val1[39] ),
    .S(net152),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03620_));
 sky130_fd_sc_hd__o22a_1 _06830_ (.A1(\top.findLeastValue.val2[39] ),
    .A2(net128),
    .B1(net119),
    .B2(_03620_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02047_));
 sky130_fd_sc_hd__mux2_1 _06831_ (.A0(\top.compVal[38] ),
    .A1(\top.findLeastValue.val1[38] ),
    .S(net152),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03621_));
 sky130_fd_sc_hd__o22a_1 _06832_ (.A1(\top.findLeastValue.val2[38] ),
    .A2(net128),
    .B1(net119),
    .B2(_03621_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02046_));
 sky130_fd_sc_hd__mux2_1 _06833_ (.A0(\top.compVal[37] ),
    .A1(\top.findLeastValue.val1[37] ),
    .S(net152),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03622_));
 sky130_fd_sc_hd__o22a_1 _06834_ (.A1(\top.findLeastValue.val2[37] ),
    .A2(net128),
    .B1(net118),
    .B2(_03622_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02045_));
 sky130_fd_sc_hd__mux2_1 _06835_ (.A0(\top.compVal[36] ),
    .A1(\top.findLeastValue.val1[36] ),
    .S(net152),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03623_));
 sky130_fd_sc_hd__o22a_1 _06836_ (.A1(\top.findLeastValue.val2[36] ),
    .A2(net128),
    .B1(net118),
    .B2(_03623_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02044_));
 sky130_fd_sc_hd__mux2_1 _06837_ (.A0(\top.compVal[35] ),
    .A1(\top.findLeastValue.val1[35] ),
    .S(net152),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03624_));
 sky130_fd_sc_hd__o22a_1 _06838_ (.A1(\top.findLeastValue.val2[35] ),
    .A2(net128),
    .B1(net118),
    .B2(_03624_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02043_));
 sky130_fd_sc_hd__mux2_1 _06839_ (.A0(\top.compVal[34] ),
    .A1(\top.findLeastValue.val1[34] ),
    .S(net152),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03625_));
 sky130_fd_sc_hd__o22a_1 _06840_ (.A1(\top.findLeastValue.val2[34] ),
    .A2(net128),
    .B1(net118),
    .B2(_03625_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02042_));
 sky130_fd_sc_hd__mux2_1 _06841_ (.A0(\top.compVal[33] ),
    .A1(\top.findLeastValue.val1[33] ),
    .S(net151),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03626_));
 sky130_fd_sc_hd__o22a_1 _06842_ (.A1(\top.findLeastValue.val2[33] ),
    .A2(net127),
    .B1(net118),
    .B2(_03626_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02041_));
 sky130_fd_sc_hd__mux2_1 _06843_ (.A0(\top.compVal[32] ),
    .A1(\top.findLeastValue.val1[32] ),
    .S(net151),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03627_));
 sky130_fd_sc_hd__o22a_1 _06844_ (.A1(\top.findLeastValue.val2[32] ),
    .A2(net127),
    .B1(net118),
    .B2(_03627_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02040_));
 sky130_fd_sc_hd__mux2_1 _06845_ (.A0(\top.compVal[31] ),
    .A1(\top.findLeastValue.val1[31] ),
    .S(net151),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03628_));
 sky130_fd_sc_hd__o22a_1 _06846_ (.A1(\top.findLeastValue.val2[31] ),
    .A2(net127),
    .B1(net118),
    .B2(_03628_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02039_));
 sky130_fd_sc_hd__mux2_1 _06847_ (.A0(\top.compVal[30] ),
    .A1(\top.findLeastValue.val1[30] ),
    .S(net151),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03629_));
 sky130_fd_sc_hd__o22a_1 _06848_ (.A1(\top.findLeastValue.val2[30] ),
    .A2(net127),
    .B1(net118),
    .B2(_03629_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02038_));
 sky130_fd_sc_hd__mux2_1 _06849_ (.A0(\top.compVal[29] ),
    .A1(\top.findLeastValue.val1[29] ),
    .S(net151),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03630_));
 sky130_fd_sc_hd__o22a_1 _06850_ (.A1(\top.findLeastValue.val2[29] ),
    .A2(net127),
    .B1(net118),
    .B2(_03630_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02037_));
 sky130_fd_sc_hd__mux2_1 _06851_ (.A0(\top.compVal[28] ),
    .A1(\top.findLeastValue.val1[28] ),
    .S(net151),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03631_));
 sky130_fd_sc_hd__o22a_1 _06852_ (.A1(\top.findLeastValue.val2[28] ),
    .A2(net127),
    .B1(net118),
    .B2(_03631_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02036_));
 sky130_fd_sc_hd__mux2_1 _06853_ (.A0(\top.compVal[27] ),
    .A1(\top.findLeastValue.val1[27] ),
    .S(net151),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03632_));
 sky130_fd_sc_hd__o22a_1 _06854_ (.A1(\top.findLeastValue.val2[27] ),
    .A2(net127),
    .B1(net117),
    .B2(_03632_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02035_));
 sky130_fd_sc_hd__mux2_1 _06855_ (.A0(\top.compVal[26] ),
    .A1(\top.findLeastValue.val1[26] ),
    .S(net150),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03633_));
 sky130_fd_sc_hd__o22a_1 _06856_ (.A1(\top.findLeastValue.val2[26] ),
    .A2(net126),
    .B1(net117),
    .B2(_03633_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02034_));
 sky130_fd_sc_hd__mux2_1 _06857_ (.A0(\top.compVal[25] ),
    .A1(\top.findLeastValue.val1[25] ),
    .S(net150),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03634_));
 sky130_fd_sc_hd__o22a_1 _06858_ (.A1(\top.findLeastValue.val2[25] ),
    .A2(net127),
    .B1(net117),
    .B2(_03634_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02033_));
 sky130_fd_sc_hd__mux2_1 _06859_ (.A0(\top.compVal[24] ),
    .A1(\top.findLeastValue.val1[24] ),
    .S(net156),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03635_));
 sky130_fd_sc_hd__o22a_1 _06860_ (.A1(\top.findLeastValue.val2[24] ),
    .A2(net132),
    .B1(net122),
    .B2(_03635_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02032_));
 sky130_fd_sc_hd__mux2_1 _06861_ (.A0(\top.compVal[23] ),
    .A1(\top.findLeastValue.val1[23] ),
    .S(net156),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03636_));
 sky130_fd_sc_hd__o22a_1 _06862_ (.A1(\top.findLeastValue.val2[23] ),
    .A2(net132),
    .B1(net117),
    .B2(_03636_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02031_));
 sky130_fd_sc_hd__mux2_1 _06863_ (.A0(\top.compVal[22] ),
    .A1(\top.findLeastValue.val1[22] ),
    .S(net156),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03637_));
 sky130_fd_sc_hd__o22a_1 _06864_ (.A1(\top.findLeastValue.val2[22] ),
    .A2(net132),
    .B1(net117),
    .B2(_03637_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02030_));
 sky130_fd_sc_hd__mux2_1 _06865_ (.A0(\top.compVal[21] ),
    .A1(\top.findLeastValue.val1[21] ),
    .S(net156),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03638_));
 sky130_fd_sc_hd__o22a_1 _06866_ (.A1(\top.findLeastValue.val2[21] ),
    .A2(net132),
    .B1(net117),
    .B2(_03638_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02029_));
 sky130_fd_sc_hd__mux2_1 _06867_ (.A0(\top.compVal[20] ),
    .A1(\top.findLeastValue.val1[20] ),
    .S(net156),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03639_));
 sky130_fd_sc_hd__o22a_1 _06868_ (.A1(\top.findLeastValue.val2[20] ),
    .A2(net132),
    .B1(net117),
    .B2(_03639_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02028_));
 sky130_fd_sc_hd__mux2_1 _06869_ (.A0(\top.compVal[19] ),
    .A1(\top.findLeastValue.val1[19] ),
    .S(net152),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03640_));
 sky130_fd_sc_hd__o22a_1 _06870_ (.A1(\top.findLeastValue.val2[19] ),
    .A2(net128),
    .B1(net117),
    .B2(_03640_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02027_));
 sky130_fd_sc_hd__mux2_1 _06871_ (.A0(\top.compVal[18] ),
    .A1(\top.findLeastValue.val1[18] ),
    .S(net155),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03641_));
 sky130_fd_sc_hd__o22a_1 _06872_ (.A1(\top.findLeastValue.val2[18] ),
    .A2(net131),
    .B1(net122),
    .B2(_03641_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02026_));
 sky130_fd_sc_hd__mux2_1 _06873_ (.A0(\top.compVal[17] ),
    .A1(\top.findLeastValue.val1[17] ),
    .S(net152),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03642_));
 sky130_fd_sc_hd__o22a_1 _06874_ (.A1(\top.findLeastValue.val2[17] ),
    .A2(net128),
    .B1(net121),
    .B2(_03642_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02025_));
 sky130_fd_sc_hd__mux2_1 _06875_ (.A0(\top.compVal[16] ),
    .A1(\top.findLeastValue.val1[16] ),
    .S(net155),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03643_));
 sky130_fd_sc_hd__o22a_1 _06876_ (.A1(\top.findLeastValue.val2[16] ),
    .A2(net128),
    .B1(net121),
    .B2(_03643_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02024_));
 sky130_fd_sc_hd__mux2_1 _06877_ (.A0(\top.compVal[15] ),
    .A1(\top.findLeastValue.val1[15] ),
    .S(net152),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03644_));
 sky130_fd_sc_hd__o22a_1 _06878_ (.A1(\top.findLeastValue.val2[15] ),
    .A2(net131),
    .B1(net122),
    .B2(_03644_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02023_));
 sky130_fd_sc_hd__mux2_1 _06879_ (.A0(\top.compVal[14] ),
    .A1(\top.findLeastValue.val1[14] ),
    .S(net154),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03645_));
 sky130_fd_sc_hd__o22a_1 _06880_ (.A1(\top.findLeastValue.val2[14] ),
    .A2(net130),
    .B1(net122),
    .B2(_03645_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02022_));
 sky130_fd_sc_hd__mux2_1 _06881_ (.A0(\top.compVal[13] ),
    .A1(\top.findLeastValue.val1[13] ),
    .S(net154),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03646_));
 sky130_fd_sc_hd__o22a_1 _06882_ (.A1(\top.findLeastValue.val2[13] ),
    .A2(net130),
    .B1(net120),
    .B2(_03646_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02021_));
 sky130_fd_sc_hd__mux2_1 _06883_ (.A0(\top.compVal[12] ),
    .A1(\top.findLeastValue.val1[12] ),
    .S(net154),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03647_));
 sky130_fd_sc_hd__o22a_1 _06884_ (.A1(\top.findLeastValue.val2[12] ),
    .A2(net130),
    .B1(net119),
    .B2(_03647_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02020_));
 sky130_fd_sc_hd__mux2_1 _06885_ (.A0(\top.compVal[11] ),
    .A1(\top.findLeastValue.val1[11] ),
    .S(net155),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03648_));
 sky130_fd_sc_hd__o22a_1 _06886_ (.A1(\top.findLeastValue.val2[11] ),
    .A2(net131),
    .B1(net120),
    .B2(_03648_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02019_));
 sky130_fd_sc_hd__mux2_1 _06887_ (.A0(\top.compVal[10] ),
    .A1(\top.findLeastValue.val1[10] ),
    .S(net154),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03649_));
 sky130_fd_sc_hd__o22a_1 _06888_ (.A1(\top.findLeastValue.val2[10] ),
    .A2(net130),
    .B1(net121),
    .B2(_03649_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02018_));
 sky130_fd_sc_hd__mux2_1 _06889_ (.A0(\top.compVal[9] ),
    .A1(\top.findLeastValue.val1[9] ),
    .S(net154),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03650_));
 sky130_fd_sc_hd__o22a_1 _06890_ (.A1(\top.findLeastValue.val2[9] ),
    .A2(net130),
    .B1(net120),
    .B2(_03650_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02017_));
 sky130_fd_sc_hd__mux2_1 _06891_ (.A0(\top.compVal[8] ),
    .A1(\top.findLeastValue.val1[8] ),
    .S(net154),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03651_));
 sky130_fd_sc_hd__o22a_1 _06892_ (.A1(\top.findLeastValue.val2[8] ),
    .A2(net130),
    .B1(net121),
    .B2(_03651_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02016_));
 sky130_fd_sc_hd__mux2_1 _06893_ (.A0(\top.compVal[7] ),
    .A1(\top.findLeastValue.val1[7] ),
    .S(net153),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03652_));
 sky130_fd_sc_hd__o22a_1 _06894_ (.A1(\top.findLeastValue.val2[7] ),
    .A2(net129),
    .B1(net120),
    .B2(_03652_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02015_));
 sky130_fd_sc_hd__mux2_1 _06895_ (.A0(\top.compVal[6] ),
    .A1(\top.findLeastValue.val1[6] ),
    .S(net153),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03653_));
 sky130_fd_sc_hd__o22a_1 _06896_ (.A1(\top.findLeastValue.val2[6] ),
    .A2(net129),
    .B1(net121),
    .B2(_03653_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02014_));
 sky130_fd_sc_hd__mux2_1 _06897_ (.A0(\top.compVal[5] ),
    .A1(\top.findLeastValue.val1[5] ),
    .S(net154),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03654_));
 sky130_fd_sc_hd__o22a_1 _06898_ (.A1(\top.findLeastValue.val2[5] ),
    .A2(net130),
    .B1(net120),
    .B2(_03654_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02013_));
 sky130_fd_sc_hd__mux2_1 _06899_ (.A0(\top.compVal[4] ),
    .A1(\top.findLeastValue.val1[4] ),
    .S(net153),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03655_));
 sky130_fd_sc_hd__o22a_1 _06900_ (.A1(\top.findLeastValue.val2[4] ),
    .A2(net129),
    .B1(net120),
    .B2(_03655_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02012_));
 sky130_fd_sc_hd__mux2_1 _06901_ (.A0(\top.compVal[3] ),
    .A1(\top.findLeastValue.val1[3] ),
    .S(net153),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03656_));
 sky130_fd_sc_hd__o22a_1 _06902_ (.A1(\top.findLeastValue.val2[3] ),
    .A2(net130),
    .B1(net120),
    .B2(_03656_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02011_));
 sky130_fd_sc_hd__mux2_1 _06903_ (.A0(\top.compVal[2] ),
    .A1(\top.findLeastValue.val1[2] ),
    .S(net153),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03657_));
 sky130_fd_sc_hd__o22a_1 _06904_ (.A1(\top.findLeastValue.val2[2] ),
    .A2(net129),
    .B1(net120),
    .B2(_03657_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02010_));
 sky130_fd_sc_hd__mux2_1 _06905_ (.A0(\top.compVal[1] ),
    .A1(\top.findLeastValue.val1[1] ),
    .S(net154),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03658_));
 sky130_fd_sc_hd__o22a_1 _06906_ (.A1(\top.findLeastValue.val2[1] ),
    .A2(net129),
    .B1(net120),
    .B2(_03658_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02009_));
 sky130_fd_sc_hd__mux2_1 _06907_ (.A0(\top.compVal[0] ),
    .A1(\top.findLeastValue.val1[0] ),
    .S(net154),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03659_));
 sky130_fd_sc_hd__o22a_1 _06908_ (.A1(\top.findLeastValue.val2[0] ),
    .A2(net130),
    .B1(net120),
    .B2(_03659_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02008_));
 sky130_fd_sc_hd__nor2_2 _06909_ (.A(net288),
    .B(net140),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03660_));
 sky130_fd_sc_hd__nand2_1 _06910_ (.A(_03394_),
    .B(net134),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03661_));
 sky130_fd_sc_hd__a21o_1 _06911_ (.A1(\top.findLeastValue.val1[46] ),
    .A2(net142),
    .B1(_03393_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02007_));
 sky130_fd_sc_hd__o22a_1 _06912_ (.A1(\top.findLeastValue.val1[45] ),
    .A2(net137),
    .B1(net113),
    .B2(net1654),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02006_));
 sky130_fd_sc_hd__o22a_1 _06913_ (.A1(\top.findLeastValue.val1[44] ),
    .A2(net136),
    .B1(net113),
    .B2(net1753),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02005_));
 sky130_fd_sc_hd__o22a_1 _06914_ (.A1(\top.findLeastValue.val1[43] ),
    .A2(net135),
    .B1(net113),
    .B2(net1730),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02004_));
 sky130_fd_sc_hd__o22a_1 _06915_ (.A1(\top.findLeastValue.val1[42] ),
    .A2(net137),
    .B1(net112),
    .B2(net1636),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02003_));
 sky130_fd_sc_hd__o22a_1 _06916_ (.A1(\top.findLeastValue.val1[41] ),
    .A2(net137),
    .B1(net112),
    .B2(\top.compVal[41] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02002_));
 sky130_fd_sc_hd__o22a_1 _06917_ (.A1(\top.findLeastValue.val1[40] ),
    .A2(net137),
    .B1(net112),
    .B2(\top.compVal[40] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02001_));
 sky130_fd_sc_hd__o22a_1 _06918_ (.A1(\top.findLeastValue.val1[39] ),
    .A2(net137),
    .B1(net112),
    .B2(net1764),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02000_));
 sky130_fd_sc_hd__o22a_1 _06919_ (.A1(\top.findLeastValue.val1[38] ),
    .A2(net137),
    .B1(net114),
    .B2(\top.compVal[38] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01999_));
 sky130_fd_sc_hd__o22a_1 _06920_ (.A1(\top.findLeastValue.val1[37] ),
    .A2(net137),
    .B1(net114),
    .B2(\top.compVal[37] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01998_));
 sky130_fd_sc_hd__o22a_1 _06921_ (.A1(\top.findLeastValue.val1[36] ),
    .A2(net137),
    .B1(net114),
    .B2(\top.compVal[36] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01997_));
 sky130_fd_sc_hd__o22a_1 _06922_ (.A1(\top.findLeastValue.val1[35] ),
    .A2(net137),
    .B1(net114),
    .B2(\top.compVal[35] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01996_));
 sky130_fd_sc_hd__o22a_1 _06923_ (.A1(\top.findLeastValue.val1[34] ),
    .A2(net133),
    .B1(net114),
    .B2(\top.compVal[34] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01995_));
 sky130_fd_sc_hd__o22a_1 _06924_ (.A1(\top.findLeastValue.val1[33] ),
    .A2(net133),
    .B1(net114),
    .B2(net1775),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01994_));
 sky130_fd_sc_hd__o22a_1 _06925_ (.A1(\top.findLeastValue.val1[32] ),
    .A2(net133),
    .B1(net114),
    .B2(\top.compVal[32] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01993_));
 sky130_fd_sc_hd__o22a_1 _06926_ (.A1(\top.findLeastValue.val1[31] ),
    .A2(net133),
    .B1(net114),
    .B2(net1762),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01992_));
 sky130_fd_sc_hd__o22a_1 _06927_ (.A1(\top.findLeastValue.val1[30] ),
    .A2(net133),
    .B1(net115),
    .B2(\top.compVal[30] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01991_));
 sky130_fd_sc_hd__o22a_1 _06928_ (.A1(\top.findLeastValue.val1[29] ),
    .A2(net133),
    .B1(net115),
    .B2(\top.compVal[29] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01990_));
 sky130_fd_sc_hd__o22a_1 _06929_ (.A1(\top.findLeastValue.val1[28] ),
    .A2(net133),
    .B1(net114),
    .B2(net1734),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01989_));
 sky130_fd_sc_hd__o22a_1 _06930_ (.A1(\top.findLeastValue.val1[27] ),
    .A2(net134),
    .B1(net115),
    .B2(\top.compVal[27] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01988_));
 sky130_fd_sc_hd__o22a_1 _06931_ (.A1(\top.findLeastValue.val1[26] ),
    .A2(net134),
    .B1(net115),
    .B2(\top.compVal[26] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01987_));
 sky130_fd_sc_hd__o22a_1 _06932_ (.A1(\top.findLeastValue.val1[25] ),
    .A2(net134),
    .B1(net115),
    .B2(net1667),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01986_));
 sky130_fd_sc_hd__o22a_1 _06933_ (.A1(\top.findLeastValue.val1[24] ),
    .A2(net134),
    .B1(net115),
    .B2(net1127),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01985_));
 sky130_fd_sc_hd__o22a_1 _06934_ (.A1(\top.findLeastValue.val1[23] ),
    .A2(net138),
    .B1(net115),
    .B2(net1776),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01984_));
 sky130_fd_sc_hd__o22a_1 _06935_ (.A1(\top.findLeastValue.val1[22] ),
    .A2(net139),
    .B1(net116),
    .B2(net1784),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01983_));
 sky130_fd_sc_hd__o22a_1 _06936_ (.A1(\top.findLeastValue.val1[21] ),
    .A2(net138),
    .B1(net116),
    .B2(net1701),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01982_));
 sky130_fd_sc_hd__o22a_1 _06937_ (.A1(\top.findLeastValue.val1[20] ),
    .A2(net138),
    .B1(net116),
    .B2(\top.compVal[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01981_));
 sky130_fd_sc_hd__o22a_1 _06938_ (.A1(\top.findLeastValue.val1[19] ),
    .A2(net138),
    .B1(net115),
    .B2(\top.compVal[19] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01980_));
 sky130_fd_sc_hd__o22a_1 _06939_ (.A1(\top.findLeastValue.val1[18] ),
    .A2(net138),
    .B1(net116),
    .B2(\top.compVal[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01979_));
 sky130_fd_sc_hd__o22a_1 _06940_ (.A1(\top.findLeastValue.val1[17] ),
    .A2(net137),
    .B1(net115),
    .B2(\top.compVal[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01978_));
 sky130_fd_sc_hd__o22a_1 _06941_ (.A1(\top.findLeastValue.val1[16] ),
    .A2(net138),
    .B1(net115),
    .B2(\top.compVal[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01977_));
 sky130_fd_sc_hd__o22a_1 _06942_ (.A1(\top.findLeastValue.val1[15] ),
    .A2(net138),
    .B1(net116),
    .B2(\top.compVal[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01976_));
 sky130_fd_sc_hd__o22a_1 _06943_ (.A1(\top.findLeastValue.val1[14] ),
    .A2(net139),
    .B1(net116),
    .B2(\top.compVal[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01975_));
 sky130_fd_sc_hd__o22a_1 _06944_ (.A1(\top.findLeastValue.val1[13] ),
    .A2(net136),
    .B1(net116),
    .B2(\top.compVal[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01974_));
 sky130_fd_sc_hd__o22a_1 _06945_ (.A1(\top.findLeastValue.val1[12] ),
    .A2(net136),
    .B1(net116),
    .B2(net1729),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01973_));
 sky130_fd_sc_hd__o22a_1 _06946_ (.A1(\top.findLeastValue.val1[11] ),
    .A2(net135),
    .B1(net113),
    .B2(net1731),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01972_));
 sky130_fd_sc_hd__o22a_1 _06947_ (.A1(\top.findLeastValue.val1[10] ),
    .A2(net136),
    .B1(net113),
    .B2(\top.compVal[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01971_));
 sky130_fd_sc_hd__o22a_1 _06948_ (.A1(\top.findLeastValue.val1[9] ),
    .A2(net136),
    .B1(net113),
    .B2(net1768),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01970_));
 sky130_fd_sc_hd__o22a_1 _06949_ (.A1(\top.findLeastValue.val1[8] ),
    .A2(net135),
    .B1(net113),
    .B2(net1687),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01969_));
 sky130_fd_sc_hd__o22a_1 _06950_ (.A1(\top.findLeastValue.val1[7] ),
    .A2(net135),
    .B1(net113),
    .B2(net1693),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01968_));
 sky130_fd_sc_hd__o22a_1 _06951_ (.A1(\top.findLeastValue.val1[6] ),
    .A2(net136),
    .B1(net113),
    .B2(net1793),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01967_));
 sky130_fd_sc_hd__o22a_1 _06952_ (.A1(\top.findLeastValue.val1[5] ),
    .A2(net135),
    .B1(net112),
    .B2(net1650),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01966_));
 sky130_fd_sc_hd__o22a_1 _06953_ (.A1(\top.findLeastValue.val1[4] ),
    .A2(net135),
    .B1(net112),
    .B2(\top.compVal[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01965_));
 sky130_fd_sc_hd__o22a_1 _06954_ (.A1(\top.findLeastValue.val1[3] ),
    .A2(net135),
    .B1(net112),
    .B2(net1698),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01964_));
 sky130_fd_sc_hd__o22a_1 _06955_ (.A1(\top.findLeastValue.val1[2] ),
    .A2(net135),
    .B1(net112),
    .B2(net1651),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01963_));
 sky130_fd_sc_hd__o22a_1 _06956_ (.A1(\top.findLeastValue.val1[1] ),
    .A2(net135),
    .B1(net112),
    .B2(net1712),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01962_));
 sky130_fd_sc_hd__o22a_1 _06957_ (.A1(\top.findLeastValue.val1[0] ),
    .A2(net135),
    .B1(net112),
    .B2(net1700),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01961_));
 sky130_fd_sc_hd__and3b_4 _06958_ (.A_N(net149),
    .B(_03609_),
    .C(net406),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03662_));
 sky130_fd_sc_hd__a21o_1 _06959_ (.A1(\top.findLeastValue.wipe_the_char_1 ),
    .A2(net149),
    .B1(_03662_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03663_));
 sky130_fd_sc_hd__a2bb2o_1 _06960_ (.A1_N(_02499_),
    .A2_N(net125),
    .B1(net123),
    .B2(_03663_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01960_));
 sky130_fd_sc_hd__a31o_1 _06961_ (.A1(net407),
    .A2(net287),
    .A3(net149),
    .B1(net142),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03664_));
 sky130_fd_sc_hd__o21a_1 _06962_ (.A1(net1711),
    .A2(net133),
    .B1(_03664_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01959_));
 sky130_fd_sc_hd__a32o_1 _06963_ (.A1(net1476),
    .A2(_02576_),
    .A3(_03395_),
    .B1(net287),
    .B2(net955),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01958_));
 sky130_fd_sc_hd__nor2_1 _06964_ (.A(net456),
    .B(net288),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03665_));
 sky130_fd_sc_hd__nand2_1 _06965_ (.A(_02562_),
    .B(net287),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03666_));
 sky130_fd_sc_hd__and2_1 _06966_ (.A(_02793_),
    .B(net287),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03667_));
 sky130_fd_sc_hd__a21oi_1 _06967_ (.A1(\top.findLeastValue.startup ),
    .A2(net459),
    .B1(net288),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03668_));
 sky130_fd_sc_hd__nand3_1 _06968_ (.A(net485),
    .B(net486),
    .C(_03088_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03669_));
 sky130_fd_sc_hd__nor2_1 _06969_ (.A(_03667_),
    .B(_03669_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03670_));
 sky130_fd_sc_hd__and2_1 _06970_ (.A(net483),
    .B(_03670_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03671_));
 sky130_fd_sc_hd__and3_1 _06971_ (.A(net482),
    .B(\top.findLeastValue.histo_index[5] ),
    .C(_03670_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03672_));
 sky130_fd_sc_hd__nor4_1 _06972_ (.A(_02501_),
    .B(_02502_),
    .C(_02503_),
    .D(_03669_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03673_));
 sky130_fd_sc_hd__a21boi_1 _06973_ (.A1(\top.findLeastValue.histo_index[7] ),
    .A2(_03672_),
    .B1_N(_03668_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03674_));
 sky130_fd_sc_hd__nor3_2 _06974_ (.A(\top.findLeastValue.startup ),
    .B(_02793_),
    .C(net288),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03675_));
 sky130_fd_sc_hd__a22o_1 _06975_ (.A1(\top.findLeastValue.histo_index[8] ),
    .A2(_03674_),
    .B1(_03675_),
    .B2(_03673_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01957_));
 sky130_fd_sc_hd__o21a_1 _06976_ (.A1(\top.findLeastValue.histo_index[7] ),
    .A2(_03672_),
    .B1(_03674_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01956_));
 sky130_fd_sc_hd__a21bo_1 _06977_ (.A1(\top.findLeastValue.histo_index[6] ),
    .A2(_03671_),
    .B1_N(_03668_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03676_));
 sky130_fd_sc_hd__o21ba_1 _06978_ (.A1(net1617),
    .A2(_03671_),
    .B1_N(_03676_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01955_));
 sky130_fd_sc_hd__a21bo_1 _06979_ (.A1(\top.findLeastValue.histo_index[5] ),
    .A2(_03670_),
    .B1_N(_03668_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03677_));
 sky130_fd_sc_hd__o21ba_1 _06980_ (.A1(net1694),
    .A2(_03670_),
    .B1_N(_03677_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01954_));
 sky130_fd_sc_hd__a21o_1 _06981_ (.A1(net486),
    .A2(_03088_),
    .B1(net484),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03678_));
 sky130_fd_sc_hd__a32o_1 _06982_ (.A1(_03669_),
    .A2(_03675_),
    .A3(_03678_),
    .B1(_03667_),
    .B2(net484),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01953_));
 sky130_fd_sc_hd__a32o_1 _06983_ (.A1(_03089_),
    .A2(_03185_),
    .A3(_03675_),
    .B1(_03667_),
    .B2(net486),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01952_));
 sky130_fd_sc_hd__a22o_1 _06984_ (.A1(\top.findLeastValue.histo_index[2] ),
    .A2(_03667_),
    .B1(_03675_),
    .B2(_03205_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01951_));
 sky130_fd_sc_hd__a32o_1 _06985_ (.A1(_02574_),
    .A2(_03087_),
    .A3(_03675_),
    .B1(_03667_),
    .B2(net487),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01950_));
 sky130_fd_sc_hd__mux2_1 _06986_ (.A0(_03667_),
    .A1(_03675_),
    .S(_02504_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01949_));
 sky130_fd_sc_hd__a2bb2o_1 _06987_ (.A1_N(_02505_),
    .A2_N(net125),
    .B1(_03660_),
    .B2(net1742),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01948_));
 sky130_fd_sc_hd__a22o_1 _06988_ (.A1(\top.cw1[6] ),
    .A2(net148),
    .B1(_03662_),
    .B2(net482),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03679_));
 sky130_fd_sc_hd__a2bb2o_1 _06989_ (.A1_N(_02506_),
    .A2_N(net125),
    .B1(net123),
    .B2(_03679_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01947_));
 sky130_fd_sc_hd__a22o_1 _06990_ (.A1(\top.cw1[5] ),
    .A2(net148),
    .B1(_03662_),
    .B2(net483),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03680_));
 sky130_fd_sc_hd__a2bb2o_1 _06991_ (.A1_N(_02507_),
    .A2_N(net125),
    .B1(net123),
    .B2(_03680_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01946_));
 sky130_fd_sc_hd__a22o_1 _06992_ (.A1(\top.cw1[4] ),
    .A2(net148),
    .B1(_03662_),
    .B2(net484),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03681_));
 sky130_fd_sc_hd__a2bb2o_1 _06993_ (.A1_N(_02508_),
    .A2_N(net125),
    .B1(net123),
    .B2(_03681_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01945_));
 sky130_fd_sc_hd__a22o_1 _06994_ (.A1(\top.cw1[3] ),
    .A2(net148),
    .B1(_03662_),
    .B2(net486),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03682_));
 sky130_fd_sc_hd__a2bb2o_1 _06995_ (.A1_N(_02509_),
    .A2_N(net125),
    .B1(net123),
    .B2(_03682_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01944_));
 sky130_fd_sc_hd__a22o_1 _06996_ (.A1(\top.cw1[2] ),
    .A2(net148),
    .B1(_03662_),
    .B2(\top.findLeastValue.histo_index[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03683_));
 sky130_fd_sc_hd__a2bb2o_1 _06997_ (.A1_N(_02510_),
    .A2_N(net125),
    .B1(net123),
    .B2(_03683_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01943_));
 sky130_fd_sc_hd__a22o_1 _06998_ (.A1(\top.cw1[1] ),
    .A2(net148),
    .B1(_03662_),
    .B2(net487),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03684_));
 sky130_fd_sc_hd__a2bb2o_1 _06999_ (.A1_N(_02511_),
    .A2_N(net126),
    .B1(net123),
    .B2(_03684_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01942_));
 sky130_fd_sc_hd__a22o_1 _07000_ (.A1(\top.cw1[0] ),
    .A2(net148),
    .B1(_03662_),
    .B2(\top.findLeastValue.histo_index[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03685_));
 sky130_fd_sc_hd__a2bb2o_1 _07001_ (.A1_N(_02512_),
    .A2_N(net126),
    .B1(net123),
    .B2(_03685_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01941_));
 sky130_fd_sc_hd__and2_1 _07002_ (.A(net1742),
    .B(net142),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01940_));
 sky130_fd_sc_hd__and3_2 _07003_ (.A(net407),
    .B(net287),
    .C(net133),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03686_));
 sky130_fd_sc_hd__a22o_1 _07004_ (.A1(net1644),
    .A2(net140),
    .B1(_03686_),
    .B2(net482),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01939_));
 sky130_fd_sc_hd__a22o_1 _07005_ (.A1(net1664),
    .A2(net140),
    .B1(_03686_),
    .B2(net483),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01938_));
 sky130_fd_sc_hd__a22o_1 _07006_ (.A1(net1779),
    .A2(net140),
    .B1(_03686_),
    .B2(net484),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01937_));
 sky130_fd_sc_hd__a22o_1 _07007_ (.A1(net1671),
    .A2(net140),
    .B1(_03686_),
    .B2(net486),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01936_));
 sky130_fd_sc_hd__a22o_1 _07008_ (.A1(net1639),
    .A2(net140),
    .B1(_03686_),
    .B2(\top.findLeastValue.histo_index[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01935_));
 sky130_fd_sc_hd__a22o_1 _07009_ (.A1(\top.cw1[1] ),
    .A2(net140),
    .B1(_03686_),
    .B2(net487),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01934_));
 sky130_fd_sc_hd__a22o_1 _07010_ (.A1(\top.cw1[0] ),
    .A2(net140),
    .B1(_03686_),
    .B2(\top.findLeastValue.histo_index[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01933_));
 sky130_fd_sc_hd__and4_1 _07011_ (.A(\top.findLeastValue.val2[10] ),
    .B(\top.findLeastValue.val2[9] ),
    .C(\top.findLeastValue.val2[8] ),
    .D(\top.findLeastValue.val2[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03687_));
 sky130_fd_sc_hd__and4_1 _07012_ (.A(\top.findLeastValue.val2[14] ),
    .B(\top.findLeastValue.val2[13] ),
    .C(\top.findLeastValue.val2[12] ),
    .D(\top.findLeastValue.val2[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03688_));
 sky130_fd_sc_hd__and4_1 _07013_ (.A(\top.findLeastValue.val2[6] ),
    .B(\top.findLeastValue.val2[5] ),
    .C(\top.findLeastValue.val2[4] ),
    .D(\top.findLeastValue.val2[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03689_));
 sky130_fd_sc_hd__and3_1 _07014_ (.A(\top.findLeastValue.val2[2] ),
    .B(\top.findLeastValue.val2[1] ),
    .C(\top.findLeastValue.val2[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03690_));
 sky130_fd_sc_hd__and4_1 _07015_ (.A(_03687_),
    .B(_03688_),
    .C(_03689_),
    .D(_03690_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03691_));
 sky130_fd_sc_hd__and4_1 _07016_ (.A(\top.findLeastValue.val2[26] ),
    .B(\top.findLeastValue.val2[25] ),
    .C(\top.findLeastValue.val2[24] ),
    .D(\top.findLeastValue.val2[23] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03692_));
 sky130_fd_sc_hd__and4_1 _07017_ (.A(\top.findLeastValue.val2[30] ),
    .B(\top.findLeastValue.val2[29] ),
    .C(\top.findLeastValue.val2[28] ),
    .D(\top.findLeastValue.val2[27] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03693_));
 sky130_fd_sc_hd__and4_1 _07018_ (.A(\top.findLeastValue.val2[22] ),
    .B(\top.findLeastValue.val2[21] ),
    .C(\top.findLeastValue.val2[20] ),
    .D(\top.findLeastValue.val2[19] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03694_));
 sky130_fd_sc_hd__and4_1 _07019_ (.A(\top.findLeastValue.val2[18] ),
    .B(\top.findLeastValue.val2[17] ),
    .C(\top.findLeastValue.val2[16] ),
    .D(\top.findLeastValue.val2[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03695_));
 sky130_fd_sc_hd__and4_1 _07020_ (.A(_03692_),
    .B(_03693_),
    .C(_03694_),
    .D(_03695_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03696_));
 sky130_fd_sc_hd__and4_1 _07021_ (.A(\top.findLeastValue.val2[42] ),
    .B(\top.findLeastValue.val2[41] ),
    .C(\top.findLeastValue.val2[40] ),
    .D(\top.findLeastValue.val2[39] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03697_));
 sky130_fd_sc_hd__and4_1 _07022_ (.A(\top.findLeastValue.val2[46] ),
    .B(\top.findLeastValue.val2[45] ),
    .C(\top.findLeastValue.val2[44] ),
    .D(\top.findLeastValue.val2[43] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03698_));
 sky130_fd_sc_hd__and4_1 _07023_ (.A(\top.findLeastValue.val2[38] ),
    .B(\top.findLeastValue.val2[37] ),
    .C(\top.findLeastValue.val2[36] ),
    .D(\top.findLeastValue.val2[35] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03699_));
 sky130_fd_sc_hd__and4_1 _07024_ (.A(\top.findLeastValue.val2[34] ),
    .B(\top.findLeastValue.val2[33] ),
    .C(\top.findLeastValue.val2[32] ),
    .D(\top.findLeastValue.val2[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03700_));
 sky130_fd_sc_hd__and4_1 _07025_ (.A(_03697_),
    .B(_03698_),
    .C(_03699_),
    .D(_03700_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03701_));
 sky130_fd_sc_hd__a31o_1 _07026_ (.A1(_03691_),
    .A2(_03696_),
    .A3(_03701_),
    .B1(_02562_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03702_));
 sky130_fd_sc_hd__and4_1 _07027_ (.A(\top.findLeastValue.val1[10] ),
    .B(\top.findLeastValue.val1[9] ),
    .C(\top.findLeastValue.val1[8] ),
    .D(\top.findLeastValue.val1[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03703_));
 sky130_fd_sc_hd__and4_1 _07028_ (.A(\top.findLeastValue.val1[14] ),
    .B(\top.findLeastValue.val1[13] ),
    .C(\top.findLeastValue.val1[12] ),
    .D(\top.findLeastValue.val1[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03704_));
 sky130_fd_sc_hd__and4_1 _07029_ (.A(\top.findLeastValue.val1[6] ),
    .B(\top.findLeastValue.val1[5] ),
    .C(\top.findLeastValue.val1[4] ),
    .D(\top.findLeastValue.val1[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03705_));
 sky130_fd_sc_hd__and3_1 _07030_ (.A(\top.findLeastValue.val1[2] ),
    .B(\top.findLeastValue.val1[1] ),
    .C(\top.findLeastValue.val1[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03706_));
 sky130_fd_sc_hd__and4_1 _07031_ (.A(_03703_),
    .B(_03704_),
    .C(_03705_),
    .D(_03706_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03707_));
 sky130_fd_sc_hd__and4_1 _07032_ (.A(\top.findLeastValue.val1[42] ),
    .B(\top.findLeastValue.val1[41] ),
    .C(\top.findLeastValue.val1[40] ),
    .D(\top.findLeastValue.val1[39] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03708_));
 sky130_fd_sc_hd__and4_1 _07033_ (.A(\top.findLeastValue.val1[46] ),
    .B(\top.findLeastValue.val1[45] ),
    .C(\top.findLeastValue.val1[44] ),
    .D(\top.findLeastValue.val1[43] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03709_));
 sky130_fd_sc_hd__and4_1 _07034_ (.A(\top.findLeastValue.val1[38] ),
    .B(\top.findLeastValue.val1[37] ),
    .C(\top.findLeastValue.val1[36] ),
    .D(\top.findLeastValue.val1[35] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03710_));
 sky130_fd_sc_hd__and4_1 _07035_ (.A(\top.findLeastValue.val1[34] ),
    .B(\top.findLeastValue.val1[33] ),
    .C(\top.findLeastValue.val1[32] ),
    .D(\top.findLeastValue.val1[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03711_));
 sky130_fd_sc_hd__and4_1 _07036_ (.A(_03708_),
    .B(_03709_),
    .C(_03710_),
    .D(_03711_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03712_));
 sky130_fd_sc_hd__and4_1 _07037_ (.A(\top.findLeastValue.val1[26] ),
    .B(\top.findLeastValue.val1[25] ),
    .C(\top.findLeastValue.val1[24] ),
    .D(\top.findLeastValue.val1[23] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03713_));
 sky130_fd_sc_hd__and4_1 _07038_ (.A(\top.findLeastValue.val1[30] ),
    .B(\top.findLeastValue.val1[29] ),
    .C(\top.findLeastValue.val1[28] ),
    .D(\top.findLeastValue.val1[27] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03714_));
 sky130_fd_sc_hd__and4_1 _07039_ (.A(\top.findLeastValue.val1[22] ),
    .B(\top.findLeastValue.val1[21] ),
    .C(\top.findLeastValue.val1[20] ),
    .D(\top.findLeastValue.val1[19] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03715_));
 sky130_fd_sc_hd__and4_1 _07040_ (.A(\top.findLeastValue.val1[18] ),
    .B(\top.findLeastValue.val1[17] ),
    .C(\top.findLeastValue.val1[16] ),
    .D(\top.findLeastValue.val1[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03716_));
 sky130_fd_sc_hd__and4_1 _07041_ (.A(_03713_),
    .B(_03714_),
    .C(_03715_),
    .D(_03716_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03717_));
 sky130_fd_sc_hd__a31o_1 _07042_ (.A1(_03707_),
    .A2(_03712_),
    .A3(_03717_),
    .B1(_03702_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03718_));
 sky130_fd_sc_hd__and2_1 _07043_ (.A(_03394_),
    .B(_03718_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03719_));
 sky130_fd_sc_hd__nor2_1 _07044_ (.A(_02455_),
    .B(_02480_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03720_));
 sky130_fd_sc_hd__xor2_1 _07045_ (.A(\top.findLeastValue.val2[39] ),
    .B(\top.findLeastValue.val1[39] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03721_));
 sky130_fd_sc_hd__nand2_1 _07046_ (.A(\top.findLeastValue.val2[38] ),
    .B(\top.findLeastValue.val1[38] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03722_));
 sky130_fd_sc_hd__or2_1 _07047_ (.A(\top.findLeastValue.val2[38] ),
    .B(\top.findLeastValue.val1[38] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03723_));
 sky130_fd_sc_hd__nand2_1 _07048_ (.A(_03722_),
    .B(_03723_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03724_));
 sky130_fd_sc_hd__nand3_1 _07049_ (.A(_03721_),
    .B(_03722_),
    .C(_03723_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03725_));
 sky130_fd_sc_hd__nor2_1 _07050_ (.A(_02460_),
    .B(_02486_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03726_));
 sky130_fd_sc_hd__nand2_1 _07051_ (.A(\top.findLeastValue.val2[37] ),
    .B(\top.findLeastValue.val1[37] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03727_));
 sky130_fd_sc_hd__nor2_1 _07052_ (.A(\top.findLeastValue.val2[37] ),
    .B(\top.findLeastValue.val1[37] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03728_));
 sky130_fd_sc_hd__nor2_1 _07053_ (.A(_03726_),
    .B(_03728_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03729_));
 sky130_fd_sc_hd__nand2_1 _07054_ (.A(\top.findLeastValue.val2[36] ),
    .B(\top.findLeastValue.val1[36] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03730_));
 sky130_fd_sc_hd__or2_1 _07055_ (.A(\top.findLeastValue.val2[36] ),
    .B(\top.findLeastValue.val1[36] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03731_));
 sky130_fd_sc_hd__nand2_1 _07056_ (.A(_03730_),
    .B(_03731_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03732_));
 sky130_fd_sc_hd__or4_2 _07057_ (.A(_03725_),
    .B(_03726_),
    .C(_03728_),
    .D(_03732_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03733_));
 sky130_fd_sc_hd__a21oi_1 _07058_ (.A1(_02459_),
    .A2(_02484_),
    .B1(_03722_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03734_));
 sky130_fd_sc_hd__a21oi_1 _07059_ (.A1(\top.findLeastValue.val2[39] ),
    .A2(\top.findLeastValue.val1[39] ),
    .B1(_03734_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03735_));
 sky130_fd_sc_hd__a211o_1 _07060_ (.A1(_03727_),
    .A2(_03730_),
    .B1(_03728_),
    .C1(_03725_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03736_));
 sky130_fd_sc_hd__nand2_1 _07061_ (.A(\top.findLeastValue.val2[24] ),
    .B(\top.findLeastValue.val1[24] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03737_));
 sky130_fd_sc_hd__a22o_1 _07062_ (.A1(\top.findLeastValue.val2[25] ),
    .A2(\top.findLeastValue.val1[25] ),
    .B1(\top.findLeastValue.val1[24] ),
    .B2(\top.findLeastValue.val2[24] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03738_));
 sky130_fd_sc_hd__o21ai_1 _07063_ (.A1(\top.findLeastValue.val2[25] ),
    .A2(\top.findLeastValue.val1[25] ),
    .B1(_03738_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03739_));
 sky130_fd_sc_hd__xor2_1 _07064_ (.A(\top.findLeastValue.val2[31] ),
    .B(\top.findLeastValue.val1[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03740_));
 sky130_fd_sc_hd__xor2_1 _07065_ (.A(\top.findLeastValue.val2[30] ),
    .B(\top.findLeastValue.val1[30] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03741_));
 sky130_fd_sc_hd__nand2_1 _07066_ (.A(_03740_),
    .B(_03741_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03742_));
 sky130_fd_sc_hd__nand2_1 _07067_ (.A(\top.findLeastValue.val2[29] ),
    .B(\top.findLeastValue.val1[29] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03743_));
 sky130_fd_sc_hd__nor2_1 _07068_ (.A(\top.findLeastValue.val2[29] ),
    .B(\top.findLeastValue.val1[29] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03744_));
 sky130_fd_sc_hd__or2_1 _07069_ (.A(\top.findLeastValue.val2[29] ),
    .B(\top.findLeastValue.val1[29] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03745_));
 sky130_fd_sc_hd__and2_1 _07070_ (.A(_03743_),
    .B(_03745_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03746_));
 sky130_fd_sc_hd__nand2_1 _07071_ (.A(\top.findLeastValue.val2[28] ),
    .B(\top.findLeastValue.val1[28] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03747_));
 sky130_fd_sc_hd__or2_1 _07072_ (.A(\top.findLeastValue.val2[28] ),
    .B(\top.findLeastValue.val1[28] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03748_));
 sky130_fd_sc_hd__nand2_1 _07073_ (.A(_03747_),
    .B(_03748_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03749_));
 sky130_fd_sc_hd__or4b_2 _07074_ (.A(_03742_),
    .B(_03749_),
    .C(_03744_),
    .D_N(_03743_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03750_));
 sky130_fd_sc_hd__nand2_1 _07075_ (.A(\top.findLeastValue.val2[26] ),
    .B(\top.findLeastValue.val1[26] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03751_));
 sky130_fd_sc_hd__or2_1 _07076_ (.A(\top.findLeastValue.val2[26] ),
    .B(\top.findLeastValue.val1[26] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03752_));
 sky130_fd_sc_hd__nand2_1 _07077_ (.A(_03751_),
    .B(_03752_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03753_));
 sky130_fd_sc_hd__nor2_1 _07078_ (.A(\top.findLeastValue.val2[27] ),
    .B(\top.findLeastValue.val1[27] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03754_));
 sky130_fd_sc_hd__and2_1 _07079_ (.A(\top.findLeastValue.val2[27] ),
    .B(\top.findLeastValue.val1[27] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03755_));
 sky130_fd_sc_hd__nor2_1 _07080_ (.A(_03754_),
    .B(_03755_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03756_));
 sky130_fd_sc_hd__or3_1 _07081_ (.A(_03753_),
    .B(_03754_),
    .C(_03755_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03757_));
 sky130_fd_sc_hd__a211oi_1 _07082_ (.A1(_03743_),
    .A2(_03747_),
    .B1(_03744_),
    .C1(_03742_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03758_));
 sky130_fd_sc_hd__o211a_1 _07083_ (.A1(\top.findLeastValue.val2[31] ),
    .A2(\top.findLeastValue.val1[31] ),
    .B1(\top.findLeastValue.val1[30] ),
    .C1(\top.findLeastValue.val2[30] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03759_));
 sky130_fd_sc_hd__a211oi_1 _07084_ (.A1(\top.findLeastValue.val2[31] ),
    .A2(\top.findLeastValue.val1[31] ),
    .B1(_03758_),
    .C1(_03759_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03760_));
 sky130_fd_sc_hd__o21ba_1 _07085_ (.A1(_03751_),
    .A2(_03754_),
    .B1_N(_03755_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03761_));
 sky130_fd_sc_hd__o21a_1 _07086_ (.A1(_03739_),
    .A2(_03757_),
    .B1(_03761_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03762_));
 sky130_fd_sc_hd__xor2_1 _07087_ (.A(\top.findLeastValue.val2[23] ),
    .B(\top.findLeastValue.val1[23] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03763_));
 sky130_fd_sc_hd__nand2_1 _07088_ (.A(\top.findLeastValue.val2[22] ),
    .B(\top.findLeastValue.val1[22] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03764_));
 sky130_fd_sc_hd__or2_1 _07089_ (.A(\top.findLeastValue.val2[22] ),
    .B(\top.findLeastValue.val1[22] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03765_));
 sky130_fd_sc_hd__nand2_1 _07090_ (.A(_03764_),
    .B(_03765_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03766_));
 sky130_fd_sc_hd__nand3_1 _07091_ (.A(_03763_),
    .B(_03764_),
    .C(_03765_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03767_));
 sky130_fd_sc_hd__xor2_2 _07092_ (.A(\top.findLeastValue.val2[18] ),
    .B(\top.findLeastValue.val1[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03768_));
 sky130_fd_sc_hd__xor2_1 _07093_ (.A(\top.findLeastValue.val2[19] ),
    .B(\top.findLeastValue.val1[19] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03769_));
 sky130_fd_sc_hd__or2_1 _07094_ (.A(\top.findLeastValue.val2[17] ),
    .B(\top.findLeastValue.val1[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03770_));
 sky130_fd_sc_hd__nand2_1 _07095_ (.A(\top.findLeastValue.val2[17] ),
    .B(\top.findLeastValue.val1[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03771_));
 sky130_fd_sc_hd__nand2_1 _07096_ (.A(\top.findLeastValue.val2[16] ),
    .B(\top.findLeastValue.val1[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03772_));
 sky130_fd_sc_hd__nand2_1 _07097_ (.A(_03771_),
    .B(_03772_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03773_));
 sky130_fd_sc_hd__and4_1 _07098_ (.A(_03768_),
    .B(_03769_),
    .C(_03770_),
    .D(_03773_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03774_));
 sky130_fd_sc_hd__o211a_1 _07099_ (.A1(\top.findLeastValue.val2[19] ),
    .A2(\top.findLeastValue.val1[19] ),
    .B1(\top.findLeastValue.val1[18] ),
    .C1(\top.findLeastValue.val2[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03775_));
 sky130_fd_sc_hd__a211o_1 _07100_ (.A1(\top.findLeastValue.val2[19] ),
    .A2(\top.findLeastValue.val1[19] ),
    .B1(_03774_),
    .C1(_03775_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03776_));
 sky130_fd_sc_hd__nand2_1 _07101_ (.A(\top.findLeastValue.val2[21] ),
    .B(\top.findLeastValue.val1[21] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03777_));
 sky130_fd_sc_hd__inv_2 _07102_ (.A(_03777_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03778_));
 sky130_fd_sc_hd__nor2_1 _07103_ (.A(\top.findLeastValue.val2[21] ),
    .B(\top.findLeastValue.val1[21] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03779_));
 sky130_fd_sc_hd__nor2_1 _07104_ (.A(_03778_),
    .B(_03779_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03780_));
 sky130_fd_sc_hd__nand2_1 _07105_ (.A(\top.findLeastValue.val2[20] ),
    .B(\top.findLeastValue.val1[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03781_));
 sky130_fd_sc_hd__or2_1 _07106_ (.A(\top.findLeastValue.val2[20] ),
    .B(\top.findLeastValue.val1[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03782_));
 sky130_fd_sc_hd__and2_1 _07107_ (.A(_03781_),
    .B(_03782_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03783_));
 sky130_fd_sc_hd__nand2_1 _07108_ (.A(_03780_),
    .B(_03783_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03784_));
 sky130_fd_sc_hd__nand2b_1 _07109_ (.A_N(_03784_),
    .B(_03776_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03785_));
 sky130_fd_sc_hd__a21o_1 _07110_ (.A1(_03777_),
    .A2(_03781_),
    .B1(_03779_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03786_));
 sky130_fd_sc_hd__a21oi_1 _07111_ (.A1(_03785_),
    .A2(_03786_),
    .B1(_03767_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03787_));
 sky130_fd_sc_hd__o211a_1 _07112_ (.A1(\top.findLeastValue.val2[23] ),
    .A2(\top.findLeastValue.val1[23] ),
    .B1(\top.findLeastValue.val1[22] ),
    .C1(\top.findLeastValue.val2[22] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03788_));
 sky130_fd_sc_hd__a211o_1 _07113_ (.A1(\top.findLeastValue.val2[23] ),
    .A2(\top.findLeastValue.val1[23] ),
    .B1(_03787_),
    .C1(_03788_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03789_));
 sky130_fd_sc_hd__nand2_1 _07114_ (.A(\top.findLeastValue.val2[14] ),
    .B(\top.findLeastValue.val1[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03790_));
 sky130_fd_sc_hd__or2_1 _07115_ (.A(\top.findLeastValue.val2[14] ),
    .B(\top.findLeastValue.val1[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03791_));
 sky130_fd_sc_hd__nand2_1 _07116_ (.A(_03790_),
    .B(_03791_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03792_));
 sky130_fd_sc_hd__nand2_1 _07117_ (.A(\top.findLeastValue.val2[15] ),
    .B(\top.findLeastValue.val1[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03793_));
 sky130_fd_sc_hd__or2_1 _07118_ (.A(\top.findLeastValue.val2[15] ),
    .B(\top.findLeastValue.val1[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03794_));
 sky130_fd_sc_hd__and2_1 _07119_ (.A(_03793_),
    .B(_03794_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03795_));
 sky130_fd_sc_hd__and3_1 _07120_ (.A(_03790_),
    .B(_03791_),
    .C(_03795_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03796_));
 sky130_fd_sc_hd__and2_1 _07121_ (.A(\top.findLeastValue.val2[12] ),
    .B(\top.findLeastValue.val1[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03797_));
 sky130_fd_sc_hd__nor2_1 _07122_ (.A(\top.findLeastValue.val2[12] ),
    .B(\top.findLeastValue.val1[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03798_));
 sky130_fd_sc_hd__nor2_1 _07123_ (.A(_03797_),
    .B(_03798_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03799_));
 sky130_fd_sc_hd__nor2_1 _07124_ (.A(_02473_),
    .B(_02495_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03800_));
 sky130_fd_sc_hd__nand2_1 _07125_ (.A(\top.findLeastValue.val2[13] ),
    .B(\top.findLeastValue.val1[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03801_));
 sky130_fd_sc_hd__or2_1 _07126_ (.A(\top.findLeastValue.val2[13] ),
    .B(\top.findLeastValue.val1[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03802_));
 sky130_fd_sc_hd__nand4_1 _07127_ (.A(_03796_),
    .B(_03799_),
    .C(_03801_),
    .D(_03802_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03803_));
 sky130_fd_sc_hd__nor2_1 _07128_ (.A(_02474_),
    .B(_02496_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03804_));
 sky130_fd_sc_hd__nor2_1 _07129_ (.A(\top.findLeastValue.val2[10] ),
    .B(\top.findLeastValue.val1[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03805_));
 sky130_fd_sc_hd__nor2_1 _07130_ (.A(_03804_),
    .B(_03805_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03806_));
 sky130_fd_sc_hd__nor2_1 _07131_ (.A(\top.findLeastValue.val2[11] ),
    .B(\top.findLeastValue.val1[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03807_));
 sky130_fd_sc_hd__or2_1 _07132_ (.A(\top.findLeastValue.val2[11] ),
    .B(\top.findLeastValue.val1[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03808_));
 sky130_fd_sc_hd__and2_1 _07133_ (.A(\top.findLeastValue.val2[11] ),
    .B(\top.findLeastValue.val1[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03809_));
 sky130_fd_sc_hd__nor2_1 _07134_ (.A(_03807_),
    .B(_03809_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03810_));
 sky130_fd_sc_hd__and2_1 _07135_ (.A(_03806_),
    .B(_03810_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03811_));
 sky130_fd_sc_hd__or2_1 _07136_ (.A(\top.findLeastValue.val2[9] ),
    .B(\top.findLeastValue.val1[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03812_));
 sky130_fd_sc_hd__nand2_1 _07137_ (.A(\top.findLeastValue.val2[9] ),
    .B(\top.findLeastValue.val1[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03813_));
 sky130_fd_sc_hd__o21ai_1 _07138_ (.A1(_02476_),
    .A2(_02497_),
    .B1(_03813_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03814_));
 sky130_fd_sc_hd__a31o_1 _07139_ (.A1(_03811_),
    .A2(_03812_),
    .A3(_03814_),
    .B1(_03809_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03815_));
 sky130_fd_sc_hd__a31o_1 _07140_ (.A1(\top.findLeastValue.val2[10] ),
    .A2(\top.findLeastValue.val1[10] ),
    .A3(_03808_),
    .B1(_03815_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03816_));
 sky130_fd_sc_hd__nor2_1 _07141_ (.A(\top.findLeastValue.val2[5] ),
    .B(\top.findLeastValue.val1[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03817_));
 sky130_fd_sc_hd__or2_1 _07142_ (.A(\top.findLeastValue.val2[5] ),
    .B(\top.findLeastValue.val1[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03818_));
 sky130_fd_sc_hd__nor2_1 _07143_ (.A(_02477_),
    .B(_02498_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03819_));
 sky130_fd_sc_hd__nand2_1 _07144_ (.A(\top.findLeastValue.val2[4] ),
    .B(\top.findLeastValue.val1[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03820_));
 sky130_fd_sc_hd__inv_2 _07145_ (.A(_03820_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03821_));
 sky130_fd_sc_hd__or2_1 _07146_ (.A(\top.findLeastValue.val2[4] ),
    .B(\top.findLeastValue.val1[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03822_));
 sky130_fd_sc_hd__and2_1 _07147_ (.A(\top.findLeastValue.val2[3] ),
    .B(\top.findLeastValue.val1[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03823_));
 sky130_fd_sc_hd__nand2_1 _07148_ (.A(\top.findLeastValue.val2[3] ),
    .B(\top.findLeastValue.val1[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03824_));
 sky130_fd_sc_hd__nand2_1 _07149_ (.A(\top.findLeastValue.val2[2] ),
    .B(\top.findLeastValue.val1[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03825_));
 sky130_fd_sc_hd__inv_2 _07150_ (.A(_03825_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03826_));
 sky130_fd_sc_hd__and2_1 _07151_ (.A(\top.findLeastValue.val2[1] ),
    .B(\top.findLeastValue.val1[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03827_));
 sky130_fd_sc_hd__xor2_1 _07152_ (.A(\top.findLeastValue.val2[1] ),
    .B(\top.findLeastValue.val1[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03828_));
 sky130_fd_sc_hd__nand2_1 _07153_ (.A(\top.findLeastValue.val2[0] ),
    .B(\top.findLeastValue.val1[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03829_));
 sky130_fd_sc_hd__and3_1 _07154_ (.A(\top.findLeastValue.val2[0] ),
    .B(\top.findLeastValue.val1[0] ),
    .C(_03828_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03830_));
 sky130_fd_sc_hd__inv_2 _07155_ (.A(_03830_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03831_));
 sky130_fd_sc_hd__or2_1 _07156_ (.A(\top.findLeastValue.val2[2] ),
    .B(\top.findLeastValue.val1[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03832_));
 sky130_fd_sc_hd__o211a_1 _07157_ (.A1(_03827_),
    .A2(_03830_),
    .B1(_03832_),
    .C1(_03825_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03833_));
 sky130_fd_sc_hd__inv_2 _07158_ (.A(_03833_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03834_));
 sky130_fd_sc_hd__or2_1 _07159_ (.A(\top.findLeastValue.val2[3] ),
    .B(\top.findLeastValue.val1[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03835_));
 sky130_fd_sc_hd__o211a_1 _07160_ (.A1(_03826_),
    .A2(_03833_),
    .B1(_03835_),
    .C1(_03824_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03836_));
 sky130_fd_sc_hd__inv_2 _07161_ (.A(_03836_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03837_));
 sky130_fd_sc_hd__o211a_1 _07162_ (.A1(_03823_),
    .A2(_03836_),
    .B1(_03820_),
    .C1(_03822_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03838_));
 sky130_fd_sc_hd__inv_2 _07163_ (.A(_03838_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03839_));
 sky130_fd_sc_hd__or2_1 _07164_ (.A(_03821_),
    .B(_03838_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03840_));
 sky130_fd_sc_hd__nor2_1 _07165_ (.A(_03817_),
    .B(_03819_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03841_));
 sky130_fd_sc_hd__o31a_1 _07166_ (.A1(_03819_),
    .A2(_03821_),
    .A3(_03838_),
    .B1(_03818_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03842_));
 sky130_fd_sc_hd__and2_1 _07167_ (.A(\top.findLeastValue.val2[7] ),
    .B(\top.findLeastValue.val1[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03843_));
 sky130_fd_sc_hd__or2_1 _07168_ (.A(\top.findLeastValue.val2[7] ),
    .B(\top.findLeastValue.val1[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03844_));
 sky130_fd_sc_hd__nand2_1 _07169_ (.A(\top.findLeastValue.val2[6] ),
    .B(\top.findLeastValue.val1[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03845_));
 sky130_fd_sc_hd__a31o_1 _07170_ (.A1(\top.findLeastValue.val2[6] ),
    .A2(\top.findLeastValue.val1[6] ),
    .A3(_03844_),
    .B1(_03843_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03846_));
 sky130_fd_sc_hd__or2_1 _07171_ (.A(\top.findLeastValue.val2[6] ),
    .B(\top.findLeastValue.val1[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03847_));
 sky130_fd_sc_hd__o221a_1 _07172_ (.A1(_03842_),
    .A2(_03846_),
    .B1(_03847_),
    .B2(_03843_),
    .C1(_03844_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03848_));
 sky130_fd_sc_hd__xor2_1 _07173_ (.A(\top.findLeastValue.val2[8] ),
    .B(\top.findLeastValue.val1[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03849_));
 sky130_fd_sc_hd__and2_1 _07174_ (.A(_03848_),
    .B(_03849_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03850_));
 sky130_fd_sc_hd__and2_1 _07175_ (.A(_03812_),
    .B(_03813_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03851_));
 sky130_fd_sc_hd__a31oi_2 _07176_ (.A1(_03811_),
    .A2(_03850_),
    .A3(_03851_),
    .B1(_03816_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03852_));
 sky130_fd_sc_hd__and2b_1 _07177_ (.A_N(_03803_),
    .B(_03816_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03853_));
 sky130_fd_sc_hd__and4b_1 _07178_ (.A_N(_03803_),
    .B(_03811_),
    .C(_03849_),
    .D(_03851_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03854_));
 sky130_fd_sc_hd__a21oi_4 _07179_ (.A1(_03848_),
    .A2(_03854_),
    .B1(_03853_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03855_));
 sky130_fd_sc_hd__a21o_1 _07180_ (.A1(_03797_),
    .A2(_03802_),
    .B1(_03800_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03856_));
 sky130_fd_sc_hd__and3_1 _07181_ (.A(\top.findLeastValue.val2[14] ),
    .B(\top.findLeastValue.val1[14] ),
    .C(_03794_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03857_));
 sky130_fd_sc_hd__a221oi_4 _07182_ (.A1(\top.findLeastValue.val2[15] ),
    .A2(\top.findLeastValue.val1[15] ),
    .B1(_03796_),
    .B2(_03856_),
    .C1(_03857_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03858_));
 sky130_fd_sc_hd__and2_1 _07183_ (.A(_03770_),
    .B(_03771_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03859_));
 sky130_fd_sc_hd__nand3_1 _07184_ (.A(_03768_),
    .B(_03769_),
    .C(_03859_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03860_));
 sky130_fd_sc_hd__or2_1 _07185_ (.A(\top.findLeastValue.val2[16] ),
    .B(\top.findLeastValue.val1[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03861_));
 sky130_fd_sc_hd__nand2_1 _07186_ (.A(_03772_),
    .B(_03861_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03862_));
 sky130_fd_sc_hd__or4_1 _07187_ (.A(_03767_),
    .B(_03784_),
    .C(_03860_),
    .D(_03862_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03863_));
 sky130_fd_sc_hd__a21oi_1 _07188_ (.A1(_03855_),
    .A2(_03858_),
    .B1(_03863_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03864_));
 sky130_fd_sc_hd__nor2_1 _07189_ (.A(_03789_),
    .B(_03864_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03865_));
 sky130_fd_sc_hd__xor2_1 _07190_ (.A(\top.findLeastValue.val2[25] ),
    .B(\top.findLeastValue.val1[25] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03866_));
 sky130_fd_sc_hd__or2_1 _07191_ (.A(\top.findLeastValue.val2[24] ),
    .B(\top.findLeastValue.val1[24] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03867_));
 sky130_fd_sc_hd__nand2_1 _07192_ (.A(_03737_),
    .B(_03867_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03868_));
 sky130_fd_sc_hd__nand3_1 _07193_ (.A(_03737_),
    .B(_03866_),
    .C(_03867_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03869_));
 sky130_fd_sc_hd__or2_1 _07194_ (.A(_03757_),
    .B(_03869_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03870_));
 sky130_fd_sc_hd__or3b_1 _07195_ (.A(_03750_),
    .B(_03870_),
    .C_N(_03789_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03871_));
 sky130_fd_sc_hd__o211a_1 _07196_ (.A1(_03750_),
    .A2(_03762_),
    .B1(_03871_),
    .C1(_03760_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03872_));
 sky130_fd_sc_hd__a2111o_1 _07197_ (.A1(_03855_),
    .A2(_03858_),
    .B1(_03863_),
    .C1(_03870_),
    .D1(_03750_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03873_));
 sky130_fd_sc_hd__and2_1 _07198_ (.A(_03872_),
    .B(_03873_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03874_));
 sky130_fd_sc_hd__nand2_1 _07199_ (.A(\top.findLeastValue.val2[34] ),
    .B(\top.findLeastValue.val1[34] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03875_));
 sky130_fd_sc_hd__or2_1 _07200_ (.A(\top.findLeastValue.val2[34] ),
    .B(\top.findLeastValue.val1[34] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03876_));
 sky130_fd_sc_hd__nand2_1 _07201_ (.A(_03875_),
    .B(_03876_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03877_));
 sky130_fd_sc_hd__nor2_1 _07202_ (.A(\top.findLeastValue.val2[35] ),
    .B(\top.findLeastValue.val1[35] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03878_));
 sky130_fd_sc_hd__nor2_1 _07203_ (.A(_02462_),
    .B(_02487_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03879_));
 sky130_fd_sc_hd__nor2_1 _07204_ (.A(_03878_),
    .B(_03879_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03880_));
 sky130_fd_sc_hd__or3_1 _07205_ (.A(_03877_),
    .B(_03878_),
    .C(_03879_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03881_));
 sky130_fd_sc_hd__nor2_1 _07206_ (.A(_02464_),
    .B(_02488_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03882_));
 sky130_fd_sc_hd__nand2_1 _07207_ (.A(\top.findLeastValue.val2[33] ),
    .B(\top.findLeastValue.val1[33] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03883_));
 sky130_fd_sc_hd__nor2_1 _07208_ (.A(\top.findLeastValue.val2[33] ),
    .B(\top.findLeastValue.val1[33] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03884_));
 sky130_fd_sc_hd__nor2_1 _07209_ (.A(_03882_),
    .B(_03884_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03885_));
 sky130_fd_sc_hd__nand2_1 _07210_ (.A(\top.findLeastValue.val2[32] ),
    .B(\top.findLeastValue.val1[32] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03886_));
 sky130_fd_sc_hd__or2_1 _07211_ (.A(\top.findLeastValue.val2[32] ),
    .B(\top.findLeastValue.val1[32] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03887_));
 sky130_fd_sc_hd__nand2_1 _07212_ (.A(_03886_),
    .B(_03887_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03888_));
 sky130_fd_sc_hd__or4_1 _07213_ (.A(_03881_),
    .B(_03882_),
    .C(_03884_),
    .D(_03888_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03889_));
 sky130_fd_sc_hd__a21o_1 _07214_ (.A1(_03872_),
    .A2(_03873_),
    .B1(_03889_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03890_));
 sky130_fd_sc_hd__a21o_1 _07215_ (.A1(_03883_),
    .A2(_03886_),
    .B1(_03884_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03891_));
 sky130_fd_sc_hd__or2_1 _07216_ (.A(_03875_),
    .B(_03878_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03892_));
 sky130_fd_sc_hd__o221a_1 _07217_ (.A1(_02462_),
    .A2(_02487_),
    .B1(_03881_),
    .B2(_03891_),
    .C1(_03892_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03893_));
 sky130_fd_sc_hd__o211a_1 _07218_ (.A1(_03733_),
    .A2(_03893_),
    .B1(_03736_),
    .C1(_03735_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03894_));
 sky130_fd_sc_hd__o21ai_4 _07219_ (.A1(_03733_),
    .A2(_03890_),
    .B1(_03894_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03895_));
 sky130_fd_sc_hd__or2_1 _07220_ (.A(\top.findLeastValue.val2[40] ),
    .B(\top.findLeastValue.val1[40] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03896_));
 sky130_fd_sc_hd__nand2_1 _07221_ (.A(\top.findLeastValue.val2[40] ),
    .B(\top.findLeastValue.val1[40] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03897_));
 sky130_fd_sc_hd__and2_1 _07222_ (.A(_03896_),
    .B(_03897_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03898_));
 sky130_fd_sc_hd__nor2_1 _07223_ (.A(\top.findLeastValue.val2[41] ),
    .B(\top.findLeastValue.val1[41] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03899_));
 sky130_fd_sc_hd__nand2_1 _07224_ (.A(\top.findLeastValue.val2[41] ),
    .B(\top.findLeastValue.val1[41] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03900_));
 sky130_fd_sc_hd__and2b_1 _07225_ (.A_N(_03899_),
    .B(_03900_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03901_));
 sky130_fd_sc_hd__nand2_1 _07226_ (.A(_03898_),
    .B(_03901_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03902_));
 sky130_fd_sc_hd__inv_2 _07227_ (.A(_03902_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03903_));
 sky130_fd_sc_hd__and2_1 _07228_ (.A(\top.findLeastValue.val2[43] ),
    .B(\top.findLeastValue.val1[43] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03904_));
 sky130_fd_sc_hd__nand2_1 _07229_ (.A(\top.findLeastValue.val2[43] ),
    .B(\top.findLeastValue.val1[43] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03905_));
 sky130_fd_sc_hd__nor2_1 _07230_ (.A(\top.findLeastValue.val2[43] ),
    .B(\top.findLeastValue.val1[43] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03906_));
 sky130_fd_sc_hd__nor2_1 _07231_ (.A(_03904_),
    .B(_03906_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03907_));
 sky130_fd_sc_hd__nand2_1 _07232_ (.A(\top.findLeastValue.val2[42] ),
    .B(\top.findLeastValue.val1[42] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03908_));
 sky130_fd_sc_hd__or2_1 _07233_ (.A(\top.findLeastValue.val2[42] ),
    .B(\top.findLeastValue.val1[42] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03909_));
 sky130_fd_sc_hd__nand2_1 _07234_ (.A(_03908_),
    .B(_03909_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03910_));
 sky130_fd_sc_hd__or3_1 _07235_ (.A(_03904_),
    .B(_03906_),
    .C(_03910_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03911_));
 sky130_fd_sc_hd__nor2_1 _07236_ (.A(_03902_),
    .B(_03911_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03912_));
 sky130_fd_sc_hd__a21o_1 _07237_ (.A1(_03897_),
    .A2(_03900_),
    .B1(_03899_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03913_));
 sky130_fd_sc_hd__o221a_1 _07238_ (.A1(_03906_),
    .A2(_03908_),
    .B1(_03911_),
    .B2(_03913_),
    .C1(_03905_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03914_));
 sky130_fd_sc_hd__a21boi_1 _07239_ (.A1(_03895_),
    .A2(_03912_),
    .B1_N(_03914_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03915_));
 sky130_fd_sc_hd__nor2_1 _07240_ (.A(\top.findLeastValue.val2[44] ),
    .B(\top.findLeastValue.val1[44] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03916_));
 sky130_fd_sc_hd__or2_1 _07241_ (.A(_03720_),
    .B(_03916_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03917_));
 sky130_fd_sc_hd__nor2_1 _07242_ (.A(_03915_),
    .B(_03917_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03918_));
 sky130_fd_sc_hd__xor2_1 _07243_ (.A(\top.findLeastValue.val2[45] ),
    .B(\top.findLeastValue.val1[45] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03919_));
 sky130_fd_sc_hd__or3_1 _07244_ (.A(_03720_),
    .B(_03918_),
    .C(_03919_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03920_));
 sky130_fd_sc_hd__o21ai_1 _07245_ (.A1(_03720_),
    .A2(_03918_),
    .B1(_03919_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03921_));
 sky130_fd_sc_hd__nor2_1 _07246_ (.A(_03393_),
    .B(_03718_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03922_));
 sky130_fd_sc_hd__a32o_1 _07247_ (.A1(_03920_),
    .A2(_03921_),
    .A3(net271),
    .B1(net277),
    .B2(net1732),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01932_));
 sky130_fd_sc_hd__a21bo_1 _07248_ (.A1(_03915_),
    .A2(_03917_),
    .B1_N(net271),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03923_));
 sky130_fd_sc_hd__a2bb2o_1 _07249_ (.A1_N(_03918_),
    .A2_N(_03923_),
    .B1(\top.findLeastValue.sum[44] ),
    .B2(net277),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01931_));
 sky130_fd_sc_hd__a21boi_2 _07250_ (.A1(_03895_),
    .A2(_03903_),
    .B1_N(_03913_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03924_));
 sky130_fd_sc_hd__o21ai_1 _07251_ (.A1(_03910_),
    .A2(_03924_),
    .B1(_03908_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03925_));
 sky130_fd_sc_hd__or2_1 _07252_ (.A(_03907_),
    .B(_03925_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03926_));
 sky130_fd_sc_hd__nand2_1 _07253_ (.A(_03907_),
    .B(_03925_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03927_));
 sky130_fd_sc_hd__a32o_1 _07254_ (.A1(net271),
    .A2(_03926_),
    .A3(_03927_),
    .B1(net277),
    .B2(net1727),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01930_));
 sky130_fd_sc_hd__xor2_2 _07255_ (.A(_03910_),
    .B(_03924_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03928_));
 sky130_fd_sc_hd__a22o_1 _07256_ (.A1(net1735),
    .A2(net278),
    .B1(net272),
    .B2(_03928_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01929_));
 sky130_fd_sc_hd__a21bo_1 _07257_ (.A1(_03895_),
    .A2(_03898_),
    .B1_N(_03897_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03929_));
 sky130_fd_sc_hd__or2_1 _07258_ (.A(_03901_),
    .B(_03929_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03930_));
 sky130_fd_sc_hd__nand2_1 _07259_ (.A(_03901_),
    .B(_03929_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03931_));
 sky130_fd_sc_hd__a32o_1 _07260_ (.A1(net271),
    .A2(_03930_),
    .A3(_03931_),
    .B1(net277),
    .B2(net1791),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01928_));
 sky130_fd_sc_hd__xor2_2 _07261_ (.A(_03895_),
    .B(_03898_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03932_));
 sky130_fd_sc_hd__a22o_1 _07262_ (.A1(\top.findLeastValue.sum[40] ),
    .A2(net278),
    .B1(net272),
    .B2(_03932_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01927_));
 sky130_fd_sc_hd__a21o_1 _07263_ (.A1(_03890_),
    .A2(_03893_),
    .B1(_03732_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03933_));
 sky130_fd_sc_hd__a31o_1 _07264_ (.A1(_03727_),
    .A2(_03730_),
    .A3(_03933_),
    .B1(_03728_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03934_));
 sky130_fd_sc_hd__o21ai_1 _07265_ (.A1(_03724_),
    .A2(_03934_),
    .B1(_03722_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03935_));
 sky130_fd_sc_hd__or2_1 _07266_ (.A(_03721_),
    .B(_03935_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03936_));
 sky130_fd_sc_hd__nand2_1 _07267_ (.A(_03721_),
    .B(_03935_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03937_));
 sky130_fd_sc_hd__a32o_1 _07268_ (.A1(net270),
    .A2(_03936_),
    .A3(_03937_),
    .B1(net276),
    .B2(net1683),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01926_));
 sky130_fd_sc_hd__nand2_1 _07269_ (.A(_03724_),
    .B(_03934_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03938_));
 sky130_fd_sc_hd__o21a_1 _07270_ (.A1(_03724_),
    .A2(_03934_),
    .B1(net270),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03939_));
 sky130_fd_sc_hd__a22o_1 _07271_ (.A1(\top.findLeastValue.sum[38] ),
    .A2(net276),
    .B1(_03938_),
    .B2(_03939_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01925_));
 sky130_fd_sc_hd__nand2_1 _07272_ (.A(_03730_),
    .B(_03933_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03940_));
 sky130_fd_sc_hd__or2_1 _07273_ (.A(_03729_),
    .B(_03940_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03941_));
 sky130_fd_sc_hd__nand2_1 _07274_ (.A(_03729_),
    .B(_03940_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03942_));
 sky130_fd_sc_hd__a32o_1 _07275_ (.A1(net270),
    .A2(_03941_),
    .A3(_03942_),
    .B1(net276),
    .B2(net1696),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01924_));
 sky130_fd_sc_hd__nand3_1 _07276_ (.A(_03732_),
    .B(_03890_),
    .C(_03893_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03943_));
 sky130_fd_sc_hd__a32o_1 _07277_ (.A1(net270),
    .A2(_03933_),
    .A3(_03943_),
    .B1(net276),
    .B2(\top.findLeastValue.sum[36] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01923_));
 sky130_fd_sc_hd__o21ai_1 _07278_ (.A1(_03874_),
    .A2(_03888_),
    .B1(_03886_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03944_));
 sky130_fd_sc_hd__o211a_1 _07279_ (.A1(_03874_),
    .A2(_03888_),
    .B1(_03886_),
    .C1(_03883_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03945_));
 sky130_fd_sc_hd__or3_1 _07280_ (.A(_03877_),
    .B(_03884_),
    .C(_03945_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03946_));
 sky130_fd_sc_hd__nand2_1 _07281_ (.A(_03875_),
    .B(_03946_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03947_));
 sky130_fd_sc_hd__or2_1 _07282_ (.A(_03880_),
    .B(_03947_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03948_));
 sky130_fd_sc_hd__nand2_1 _07283_ (.A(_03880_),
    .B(_03947_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03949_));
 sky130_fd_sc_hd__a32o_1 _07284_ (.A1(net270),
    .A2(_03948_),
    .A3(_03949_),
    .B1(net276),
    .B2(\top.findLeastValue.sum[35] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01922_));
 sky130_fd_sc_hd__o21ai_1 _07285_ (.A1(_03884_),
    .A2(_03945_),
    .B1(_03877_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03950_));
 sky130_fd_sc_hd__a32o_1 _07286_ (.A1(net270),
    .A2(_03946_),
    .A3(_03950_),
    .B1(net276),
    .B2(\top.findLeastValue.sum[34] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01921_));
 sky130_fd_sc_hd__or2_1 _07287_ (.A(_03885_),
    .B(_03944_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03951_));
 sky130_fd_sc_hd__nand2_1 _07288_ (.A(_03885_),
    .B(_03944_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03952_));
 sky130_fd_sc_hd__a32o_1 _07289_ (.A1(net270),
    .A2(_03951_),
    .A3(_03952_),
    .B1(net276),
    .B2(net1715),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01920_));
 sky130_fd_sc_hd__nand2_1 _07290_ (.A(_03874_),
    .B(_03888_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03953_));
 sky130_fd_sc_hd__o21a_1 _07291_ (.A1(_03874_),
    .A2(_03888_),
    .B1(net270),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03954_));
 sky130_fd_sc_hd__a22o_1 _07292_ (.A1(\top.findLeastValue.sum[32] ),
    .A2(net276),
    .B1(_03953_),
    .B2(_03954_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01919_));
 sky130_fd_sc_hd__or2_1 _07293_ (.A(_03865_),
    .B(_03868_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03955_));
 sky130_fd_sc_hd__o21ai_1 _07294_ (.A1(_03865_),
    .A2(_03869_),
    .B1(_03739_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03956_));
 sky130_fd_sc_hd__o21bai_1 _07295_ (.A1(_03789_),
    .A2(_03864_),
    .B1_N(_03870_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03957_));
 sky130_fd_sc_hd__a21o_1 _07296_ (.A1(_03762_),
    .A2(_03957_),
    .B1(_03749_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03958_));
 sky130_fd_sc_hd__nand3_1 _07297_ (.A(_03743_),
    .B(_03747_),
    .C(_03958_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03959_));
 sky130_fd_sc_hd__nand2_1 _07298_ (.A(_03745_),
    .B(_03959_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03960_));
 sky130_fd_sc_hd__a32o_1 _07299_ (.A1(_03741_),
    .A2(_03745_),
    .A3(_03959_),
    .B1(\top.findLeastValue.val1[30] ),
    .B2(\top.findLeastValue.val2[30] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03961_));
 sky130_fd_sc_hd__or2_1 _07300_ (.A(_03740_),
    .B(_03961_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03962_));
 sky130_fd_sc_hd__nand2_1 _07301_ (.A(_03740_),
    .B(_03961_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03963_));
 sky130_fd_sc_hd__a32o_1 _07302_ (.A1(net268),
    .A2(_03962_),
    .A3(_03963_),
    .B1(net274),
    .B2(net1705),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01918_));
 sky130_fd_sc_hd__xnor2_1 _07303_ (.A(_03741_),
    .B(_03960_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03964_));
 sky130_fd_sc_hd__a22o_1 _07304_ (.A1(net1725),
    .A2(net274),
    .B1(net268),
    .B2(_03964_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01917_));
 sky130_fd_sc_hd__nand2_1 _07305_ (.A(_03747_),
    .B(_03958_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03965_));
 sky130_fd_sc_hd__or2_1 _07306_ (.A(_03746_),
    .B(_03965_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03966_));
 sky130_fd_sc_hd__nand2_1 _07307_ (.A(_03746_),
    .B(_03965_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03967_));
 sky130_fd_sc_hd__a32o_1 _07308_ (.A1(net268),
    .A2(_03966_),
    .A3(_03967_),
    .B1(net274),
    .B2(net1656),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01916_));
 sky130_fd_sc_hd__nand3_1 _07309_ (.A(_03749_),
    .B(_03762_),
    .C(_03957_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03968_));
 sky130_fd_sc_hd__a32o_1 _07310_ (.A1(net268),
    .A2(_03958_),
    .A3(_03968_),
    .B1(net274),
    .B2(net1659),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01915_));
 sky130_fd_sc_hd__a21bo_1 _07311_ (.A1(_03752_),
    .A2(_03956_),
    .B1_N(_03751_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03969_));
 sky130_fd_sc_hd__or2_1 _07312_ (.A(_03756_),
    .B(_03969_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03970_));
 sky130_fd_sc_hd__nand2_1 _07313_ (.A(_03756_),
    .B(_03969_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03971_));
 sky130_fd_sc_hd__a32o_1 _07314_ (.A1(net268),
    .A2(_03970_),
    .A3(_03971_),
    .B1(net274),
    .B2(net1676),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01914_));
 sky130_fd_sc_hd__xnor2_1 _07315_ (.A(_03753_),
    .B(_03956_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03972_));
 sky130_fd_sc_hd__a22o_1 _07316_ (.A1(net1648),
    .A2(net274),
    .B1(net268),
    .B2(_03972_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01913_));
 sky130_fd_sc_hd__nand2_1 _07317_ (.A(_03737_),
    .B(_03955_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03973_));
 sky130_fd_sc_hd__or2_1 _07318_ (.A(_03866_),
    .B(_03973_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03974_));
 sky130_fd_sc_hd__nand2_1 _07319_ (.A(_03866_),
    .B(_03973_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03975_));
 sky130_fd_sc_hd__a32o_1 _07320_ (.A1(net268),
    .A2(_03974_),
    .A3(_03975_),
    .B1(net274),
    .B2(net1669),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01912_));
 sky130_fd_sc_hd__nand2_1 _07321_ (.A(_03865_),
    .B(_03868_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03976_));
 sky130_fd_sc_hd__a32o_1 _07322_ (.A1(net268),
    .A2(_03955_),
    .A3(_03976_),
    .B1(net274),
    .B2(net1627),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01911_));
 sky130_fd_sc_hd__a21o_1 _07323_ (.A1(_03855_),
    .A2(_03858_),
    .B1(_03862_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03977_));
 sky130_fd_sc_hd__nor2_1 _07324_ (.A(_03860_),
    .B(_03977_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03978_));
 sky130_fd_sc_hd__o21ai_1 _07325_ (.A1(_03776_),
    .A2(_03978_),
    .B1(_03783_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03979_));
 sky130_fd_sc_hd__o21a_1 _07326_ (.A1(_03779_),
    .A2(_03979_),
    .B1(_03786_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03980_));
 sky130_fd_sc_hd__o21ai_1 _07327_ (.A1(_03766_),
    .A2(_03980_),
    .B1(_03764_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03981_));
 sky130_fd_sc_hd__or2_1 _07328_ (.A(_03763_),
    .B(_03981_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03982_));
 sky130_fd_sc_hd__nand2_1 _07329_ (.A(_03763_),
    .B(_03981_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03983_));
 sky130_fd_sc_hd__a32o_1 _07330_ (.A1(net268),
    .A2(_03982_),
    .A3(_03983_),
    .B1(net274),
    .B2(net1616),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01910_));
 sky130_fd_sc_hd__xor2_1 _07331_ (.A(_03766_),
    .B(_03980_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03984_));
 sky130_fd_sc_hd__a22o_1 _07332_ (.A1(net1733),
    .A2(net275),
    .B1(net269),
    .B2(_03984_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01909_));
 sky130_fd_sc_hd__nand2_1 _07333_ (.A(_03781_),
    .B(_03979_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03985_));
 sky130_fd_sc_hd__or2_1 _07334_ (.A(_03780_),
    .B(_03985_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03986_));
 sky130_fd_sc_hd__nand2_1 _07335_ (.A(_03780_),
    .B(_03985_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03987_));
 sky130_fd_sc_hd__a32o_1 _07336_ (.A1(net269),
    .A2(_03986_),
    .A3(_03987_),
    .B1(net275),
    .B2(net1680),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01908_));
 sky130_fd_sc_hd__or3_1 _07337_ (.A(_03776_),
    .B(_03783_),
    .C(_03978_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03988_));
 sky130_fd_sc_hd__a32o_1 _07338_ (.A1(net269),
    .A2(_03979_),
    .A3(_03988_),
    .B1(net275),
    .B2(net1624),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01907_));
 sky130_fd_sc_hd__nand2b_1 _07339_ (.A_N(_03773_),
    .B(_03977_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03989_));
 sky130_fd_sc_hd__nand2_1 _07340_ (.A(_03770_),
    .B(_03989_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03990_));
 sky130_fd_sc_hd__a32o_1 _07341_ (.A1(_03768_),
    .A2(_03770_),
    .A3(_03989_),
    .B1(\top.findLeastValue.val1[18] ),
    .B2(\top.findLeastValue.val2[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03991_));
 sky130_fd_sc_hd__or2_1 _07342_ (.A(_03769_),
    .B(_03991_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03992_));
 sky130_fd_sc_hd__nand2_1 _07343_ (.A(_03769_),
    .B(_03991_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03993_));
 sky130_fd_sc_hd__a32o_1 _07344_ (.A1(net268),
    .A2(_03992_),
    .A3(_03993_),
    .B1(net275),
    .B2(net1630),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01906_));
 sky130_fd_sc_hd__xnor2_1 _07345_ (.A(_03768_),
    .B(_03990_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03994_));
 sky130_fd_sc_hd__a22o_1 _07346_ (.A1(net1706),
    .A2(net274),
    .B1(net269),
    .B2(_03994_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01905_));
 sky130_fd_sc_hd__nand2_1 _07347_ (.A(_03772_),
    .B(_03977_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03995_));
 sky130_fd_sc_hd__or2_1 _07348_ (.A(_03859_),
    .B(_03995_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03996_));
 sky130_fd_sc_hd__nand2_1 _07349_ (.A(_03859_),
    .B(_03995_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03997_));
 sky130_fd_sc_hd__a32o_1 _07350_ (.A1(net269),
    .A2(_03996_),
    .A3(_03997_),
    .B1(net275),
    .B2(net1709),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01904_));
 sky130_fd_sc_hd__nand3_1 _07351_ (.A(_03855_),
    .B(_03858_),
    .C(_03862_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03998_));
 sky130_fd_sc_hd__a32o_1 _07352_ (.A1(net269),
    .A2(_03977_),
    .A3(_03998_),
    .B1(net275),
    .B2(net1707),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01903_));
 sky130_fd_sc_hd__o21bai_1 _07353_ (.A1(_03798_),
    .A2(_03852_),
    .B1_N(_03797_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_03999_));
 sky130_fd_sc_hd__a21o_1 _07354_ (.A1(_03802_),
    .A2(_03999_),
    .B1(_03800_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04000_));
 sky130_fd_sc_hd__a21bo_1 _07355_ (.A1(_03791_),
    .A2(_04000_),
    .B1_N(_03790_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04001_));
 sky130_fd_sc_hd__or2_1 _07356_ (.A(_03795_),
    .B(_04001_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04002_));
 sky130_fd_sc_hd__nand2_1 _07357_ (.A(_03795_),
    .B(_04001_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04003_));
 sky130_fd_sc_hd__a32o_1 _07358_ (.A1(net272),
    .A2(_04002_),
    .A3(_04003_),
    .B1(net278),
    .B2(\top.findLeastValue.sum[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01902_));
 sky130_fd_sc_hd__xnor2_1 _07359_ (.A(_03792_),
    .B(_04000_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04004_));
 sky130_fd_sc_hd__a22o_1 _07360_ (.A1(\top.findLeastValue.sum[14] ),
    .A2(net278),
    .B1(net272),
    .B2(_04004_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01901_));
 sky130_fd_sc_hd__a21o_1 _07361_ (.A1(_03801_),
    .A2(_03802_),
    .B1(_03999_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04005_));
 sky130_fd_sc_hd__nand3_1 _07362_ (.A(_03801_),
    .B(_03802_),
    .C(_03999_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04006_));
 sky130_fd_sc_hd__a32o_1 _07363_ (.A1(net273),
    .A2(_04005_),
    .A3(_04006_),
    .B1(net279),
    .B2(net1559),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01900_));
 sky130_fd_sc_hd__xnor2_1 _07364_ (.A(_03799_),
    .B(_03852_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04007_));
 sky130_fd_sc_hd__a22o_1 _07365_ (.A1(\top.findLeastValue.sum[12] ),
    .A2(net279),
    .B1(net272),
    .B2(_04007_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01899_));
 sky130_fd_sc_hd__o21a_1 _07366_ (.A1(_03814_),
    .A2(_03850_),
    .B1(_03812_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04008_));
 sky130_fd_sc_hd__a21o_1 _07367_ (.A1(_03806_),
    .A2(_04008_),
    .B1(_03804_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04009_));
 sky130_fd_sc_hd__or2_1 _07368_ (.A(_03810_),
    .B(_04009_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04010_));
 sky130_fd_sc_hd__nand2_1 _07369_ (.A(_03810_),
    .B(_04009_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04011_));
 sky130_fd_sc_hd__a32o_1 _07370_ (.A1(net272),
    .A2(_04010_),
    .A3(_04011_),
    .B1(net278),
    .B2(\top.findLeastValue.sum[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01898_));
 sky130_fd_sc_hd__xor2_1 _07371_ (.A(_03806_),
    .B(_04008_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04012_));
 sky130_fd_sc_hd__a22o_1 _07372_ (.A1(\top.findLeastValue.sum[10] ),
    .A2(net278),
    .B1(net272),
    .B2(_04012_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01897_));
 sky130_fd_sc_hd__a21o_1 _07373_ (.A1(\top.findLeastValue.val2[8] ),
    .A2(\top.findLeastValue.val1[8] ),
    .B1(_03850_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04013_));
 sky130_fd_sc_hd__or2_1 _07374_ (.A(_03851_),
    .B(_04013_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04014_));
 sky130_fd_sc_hd__nand2_1 _07375_ (.A(_03851_),
    .B(_04013_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04015_));
 sky130_fd_sc_hd__a32o_1 _07376_ (.A1(net273),
    .A2(_04014_),
    .A3(_04015_),
    .B1(net279),
    .B2(\top.findLeastValue.sum[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01896_));
 sky130_fd_sc_hd__or2_1 _07377_ (.A(_03848_),
    .B(_03849_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04016_));
 sky130_fd_sc_hd__and3b_1 _07378_ (.A_N(_03850_),
    .B(net273),
    .C(_04016_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04017_));
 sky130_fd_sc_hd__a21o_1 _07379_ (.A1(net1743),
    .A2(net278),
    .B1(_04017_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01895_));
 sky130_fd_sc_hd__nand3_1 _07380_ (.A(_03842_),
    .B(_03845_),
    .C(_03847_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04018_));
 sky130_fd_sc_hd__nand2_1 _07381_ (.A(_03845_),
    .B(_04018_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04019_));
 sky130_fd_sc_hd__nand2b_1 _07382_ (.A_N(_03843_),
    .B(_03844_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04020_));
 sky130_fd_sc_hd__xnor2_1 _07383_ (.A(_04019_),
    .B(_04020_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04021_));
 sky130_fd_sc_hd__a22o_1 _07384_ (.A1(net1789),
    .A2(net277),
    .B1(net272),
    .B2(_04021_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01894_));
 sky130_fd_sc_hd__a21o_1 _07385_ (.A1(_03845_),
    .A2(_03847_),
    .B1(_03842_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04022_));
 sky130_fd_sc_hd__a32o_1 _07386_ (.A1(net271),
    .A2(_04018_),
    .A3(_04022_),
    .B1(net278),
    .B2(\top.findLeastValue.sum[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01893_));
 sky130_fd_sc_hd__nand2_1 _07387_ (.A(_03840_),
    .B(_03841_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04023_));
 sky130_fd_sc_hd__or2_1 _07388_ (.A(_03840_),
    .B(_03841_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04024_));
 sky130_fd_sc_hd__a32o_1 _07389_ (.A1(net272),
    .A2(_04023_),
    .A3(_04024_),
    .B1(net278),
    .B2(\top.findLeastValue.sum[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01892_));
 sky130_fd_sc_hd__a211o_1 _07390_ (.A1(_03820_),
    .A2(_03822_),
    .B1(_03823_),
    .C1(_03836_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04025_));
 sky130_fd_sc_hd__a32o_1 _07391_ (.A1(_03839_),
    .A2(net271),
    .A3(_04025_),
    .B1(net277),
    .B2(\top.findLeastValue.sum[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01891_));
 sky130_fd_sc_hd__a211o_1 _07392_ (.A1(_03824_),
    .A2(_03835_),
    .B1(_03833_),
    .C1(_03826_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04026_));
 sky130_fd_sc_hd__a32o_1 _07393_ (.A1(_03837_),
    .A2(net271),
    .A3(_04026_),
    .B1(net277),
    .B2(\top.findLeastValue.sum[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01890_));
 sky130_fd_sc_hd__a211o_1 _07394_ (.A1(_03825_),
    .A2(_03832_),
    .B1(_03830_),
    .C1(_03827_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04027_));
 sky130_fd_sc_hd__a32o_1 _07395_ (.A1(_03834_),
    .A2(net271),
    .A3(_04027_),
    .B1(net277),
    .B2(\top.findLeastValue.sum[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01889_));
 sky130_fd_sc_hd__nand2b_1 _07396_ (.A_N(_03828_),
    .B(_03829_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04028_));
 sky130_fd_sc_hd__a32o_1 _07397_ (.A1(_03831_),
    .A2(net271),
    .A3(_04028_),
    .B1(net277),
    .B2(net1749),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01888_));
 sky130_fd_sc_hd__or2_1 _07398_ (.A(\top.findLeastValue.val2[0] ),
    .B(\top.findLeastValue.val1[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04029_));
 sky130_fd_sc_hd__a32o_1 _07399_ (.A1(_03829_),
    .A2(net271),
    .A3(_04029_),
    .B1(net277),
    .B2(net1724),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01887_));
 sky130_fd_sc_hd__a21oi_1 _07400_ (.A1(_02522_),
    .A2(net150),
    .B1(_03662_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04030_));
 sky130_fd_sc_hd__o22a_1 _07401_ (.A1(\top.findLeastValue.least2[8] ),
    .A2(_03611_),
    .B1(net117),
    .B2(_04030_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01886_));
 sky130_fd_sc_hd__mux2_1 _07402_ (.A0(\top.findLeastValue.histo_index[7] ),
    .A1(_02523_),
    .S(net148),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04031_));
 sky130_fd_sc_hd__nor2_1 _07403_ (.A(_03662_),
    .B(_04031_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04032_));
 sky130_fd_sc_hd__o22a_1 _07404_ (.A1(\top.findLeastValue.least2[7] ),
    .A2(net127),
    .B1(net117),
    .B2(_04032_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01885_));
 sky130_fd_sc_hd__mux2_1 _07405_ (.A0(net482),
    .A1(\top.findLeastValue.least1[6] ),
    .S(net150),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04033_));
 sky130_fd_sc_hd__a2bb2o_1 _07406_ (.A1_N(_02515_),
    .A2_N(net126),
    .B1(net123),
    .B2(_04033_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01884_));
 sky130_fd_sc_hd__mux2_1 _07407_ (.A0(net483),
    .A1(\top.findLeastValue.least1[5] ),
    .S(net149),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04034_));
 sky130_fd_sc_hd__a2bb2o_1 _07408_ (.A1_N(_02516_),
    .A2_N(net125),
    .B1(net124),
    .B2(_04034_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01883_));
 sky130_fd_sc_hd__mux2_1 _07409_ (.A0(net485),
    .A1(\top.findLeastValue.least1[4] ),
    .S(net150),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04035_));
 sky130_fd_sc_hd__a2bb2o_1 _07410_ (.A1_N(_02517_),
    .A2_N(net126),
    .B1(net124),
    .B2(_04035_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01882_));
 sky130_fd_sc_hd__mux2_1 _07411_ (.A0(\top.findLeastValue.histo_index[3] ),
    .A1(\top.findLeastValue.least1[3] ),
    .S(net150),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04036_));
 sky130_fd_sc_hd__a2bb2o_1 _07412_ (.A1_N(_02518_),
    .A2_N(net126),
    .B1(net124),
    .B2(_04036_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01881_));
 sky130_fd_sc_hd__mux2_1 _07413_ (.A0(\top.findLeastValue.histo_index[2] ),
    .A1(\top.findLeastValue.least1[2] ),
    .S(net148),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04037_));
 sky130_fd_sc_hd__a2bb2o_1 _07414_ (.A1_N(_02519_),
    .A2_N(net126),
    .B1(net124),
    .B2(_04037_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01880_));
 sky130_fd_sc_hd__mux2_1 _07415_ (.A0(net487),
    .A1(\top.findLeastValue.least1[1] ),
    .S(net149),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04038_));
 sky130_fd_sc_hd__a2bb2o_1 _07416_ (.A1_N(_02520_),
    .A2_N(net126),
    .B1(net124),
    .B2(_04038_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01879_));
 sky130_fd_sc_hd__mux2_1 _07417_ (.A0(\top.findLeastValue.histo_index[0] ),
    .A1(\top.findLeastValue.least1[0] ),
    .S(net148),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04039_));
 sky130_fd_sc_hd__a2bb2o_1 _07418_ (.A1_N(_02521_),
    .A2_N(net125),
    .B1(net123),
    .B2(_04039_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01878_));
 sky130_fd_sc_hd__o21ai_1 _07419_ (.A1(_02522_),
    .A2(net133),
    .B1(_03664_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_01877_));
 sky130_fd_sc_hd__a21o_1 _07420_ (.A1(_03412_),
    .A2(net149),
    .B1(_02523_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04040_));
 sky130_fd_sc_hd__nand2_1 _07421_ (.A(net287),
    .B(_04040_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_01876_));
 sky130_fd_sc_hd__a22o_1 _07422_ (.A1(\top.findLeastValue.least1[6] ),
    .A2(net141),
    .B1(_03660_),
    .B2(net482),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01875_));
 sky130_fd_sc_hd__a22o_1 _07423_ (.A1(\top.findLeastValue.least1[5] ),
    .A2(net141),
    .B1(_03660_),
    .B2(net483),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01874_));
 sky130_fd_sc_hd__a22o_1 _07424_ (.A1(\top.findLeastValue.least1[4] ),
    .A2(net141),
    .B1(_03660_),
    .B2(net485),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01873_));
 sky130_fd_sc_hd__a22o_1 _07425_ (.A1(\top.findLeastValue.least1[3] ),
    .A2(net141),
    .B1(_03660_),
    .B2(net1615),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01872_));
 sky130_fd_sc_hd__a22o_1 _07426_ (.A1(\top.findLeastValue.least1[2] ),
    .A2(net141),
    .B1(_03660_),
    .B2(\top.findLeastValue.histo_index[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01871_));
 sky130_fd_sc_hd__a22o_1 _07427_ (.A1(\top.findLeastValue.least1[1] ),
    .A2(net140),
    .B1(_03660_),
    .B2(net1143),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01870_));
 sky130_fd_sc_hd__a22o_1 _07428_ (.A1(\top.findLeastValue.least1[0] ),
    .A2(net140),
    .B1(_03660_),
    .B2(\top.findLeastValue.histo_index[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01869_));
 sky130_fd_sc_hd__o31a_1 _07429_ (.A1(\top.dut.bits_in_buf[1] ),
    .A2(\top.dut.bits_in_buf[0] ),
    .A3(\top.dut.bits_in_buf[2] ),
    .B1(net713),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04041_));
 sky130_fd_sc_hd__xnor2_1 _07430_ (.A(\top.dut.bits_in_buf[3] ),
    .B(_04041_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04042_));
 sky130_fd_sc_hd__inv_2 _07431_ (.A(net344),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\top.dut.out_valid_next ));
 sky130_fd_sc_hd__or3_2 _07432_ (.A(_02405_),
    .B(\top.dut.bits_in_buf[1] ),
    .C(\top.dut.bits_in_buf[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04043_));
 sky130_fd_sc_hd__xor2_4 _07433_ (.A(\top.dut.bits_in_buf[2] ),
    .B(_04043_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04044_));
 sky130_fd_sc_hd__inv_2 _07434_ (.A(_04044_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\top.dut.bits_in_buf_next[2] ));
 sky130_fd_sc_hd__nor2_2 _07435_ (.A(net344),
    .B(\top.dut.bits_in_buf_next[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04045_));
 sky130_fd_sc_hd__nand2_2 _07436_ (.A(\top.dut.out_valid_next ),
    .B(_04044_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04046_));
 sky130_fd_sc_hd__o21ai_1 _07437_ (.A1(_02405_),
    .A2(\top.dut.bits_in_buf[0] ),
    .B1(\top.dut.bits_in_buf[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04047_));
 sky130_fd_sc_hd__and2_1 _07438_ (.A(_04043_),
    .B(_04047_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04048_));
 sky130_fd_sc_hd__inv_2 _07439_ (.A(net342),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\top.dut.bits_in_buf_next[1] ));
 sky130_fd_sc_hd__xnor2_2 _07440_ (.A(net714),
    .B(\top.dut.bits_in_buf[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04049_));
 sky130_fd_sc_hd__inv_2 _07441_ (.A(net393),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\top.dut.bits_in_buf_next[0] ));
 sky130_fd_sc_hd__mux2_1 _07442_ (.A0(\top.dut.bit_buf[10] ),
    .A1(\top.dut.bit_buf[3] ),
    .S(net714),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04050_));
 sky130_fd_sc_hd__mux2_1 _07443_ (.A0(\top.dut.bit_buf[9] ),
    .A1(\top.dut.bit_buf[2] ),
    .S(net713),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04051_));
 sky130_fd_sc_hd__mux2_1 _07444_ (.A0(_04050_),
    .A1(_04051_),
    .S(net393),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04052_));
 sky130_fd_sc_hd__mux2_1 _07445_ (.A0(\top.dut.bit_buf[8] ),
    .A1(\top.dut.bit_buf[1] ),
    .S(net714),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04053_));
 sky130_fd_sc_hd__mux2_1 _07446_ (.A0(\top.dut.bit_buf[7] ),
    .A1(\top.dut.bit_buf[0] ),
    .S(net713),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04054_));
 sky130_fd_sc_hd__mux2_1 _07447_ (.A0(_04053_),
    .A1(_04054_),
    .S(_04049_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04055_));
 sky130_fd_sc_hd__mux2_1 _07448_ (.A0(_04052_),
    .A1(_04055_),
    .S(net342),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04056_));
 sky130_fd_sc_hd__and3_1 _07449_ (.A(\top.dut.bits_in_buf[1] ),
    .B(\top.dut.bits_in_buf[2] ),
    .C(net393),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04057_));
 sky130_fd_sc_hd__mux2_1 _07450_ (.A0(\top.dut.bit_buf[13] ),
    .A1(\top.dut.bit_buf[6] ),
    .S(net713),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04058_));
 sky130_fd_sc_hd__and2_1 _07451_ (.A(\top.dut.out[7] ),
    .B(net343),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04059_));
 sky130_fd_sc_hd__nor2_2 _07452_ (.A(net343),
    .B(_04044_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04060_));
 sky130_fd_sc_hd__or2_1 _07453_ (.A(net344),
    .B(_04044_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04061_));
 sky130_fd_sc_hd__mux2_1 _07454_ (.A0(\top.dut.bit_buf[12] ),
    .A1(\top.dut.bit_buf[5] ),
    .S(net713),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04062_));
 sky130_fd_sc_hd__mux2_1 _07455_ (.A0(\top.dut.bit_buf[11] ),
    .A1(\top.dut.bit_buf[4] ),
    .S(net713),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04063_));
 sky130_fd_sc_hd__mux2_1 _07456_ (.A0(_04062_),
    .A1(_04063_),
    .S(net393),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04064_));
 sky130_fd_sc_hd__and3_1 _07457_ (.A(_04048_),
    .B(_04060_),
    .C(_04064_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04065_));
 sky130_fd_sc_hd__a311o_1 _07458_ (.A1(\top.dut.out_valid_next ),
    .A2(_04057_),
    .A3(_04058_),
    .B1(_04059_),
    .C1(_04065_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04066_));
 sky130_fd_sc_hd__a21o_1 _07459_ (.A1(_04045_),
    .A2(_04056_),
    .B1(_04066_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01868_));
 sky130_fd_sc_hd__nor2_1 _07460_ (.A(net342),
    .B(net393),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04067_));
 sky130_fd_sc_hd__and3_1 _07461_ (.A(\top.dut.bits_in_buf[1] ),
    .B(net393),
    .C(_04062_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04068_));
 sky130_fd_sc_hd__mux2_1 _07462_ (.A0(_04050_),
    .A1(_04063_),
    .S(\top.dut.bits_in_buf_next[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04069_));
 sky130_fd_sc_hd__a221o_1 _07463_ (.A1(_04058_),
    .A2(_04067_),
    .B1(_04069_),
    .B2(_04048_),
    .C1(_04068_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04070_));
 sky130_fd_sc_hd__mux2_1 _07464_ (.A0(_04051_),
    .A1(_04053_),
    .S(net393),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04071_));
 sky130_fd_sc_hd__mux2_1 _07465_ (.A0(\top.dut.bit_buf[6] ),
    .A1(net35),
    .S(net713),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04072_));
 sky130_fd_sc_hd__mux2_1 _07466_ (.A0(_04054_),
    .A1(_04072_),
    .S(_04049_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04073_));
 sky130_fd_sc_hd__mux2_1 _07467_ (.A0(_04071_),
    .A1(_04073_),
    .S(net342),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04074_));
 sky130_fd_sc_hd__a22o_1 _07468_ (.A1(_04060_),
    .A2(_04070_),
    .B1(_04074_),
    .B2(_04045_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04075_));
 sky130_fd_sc_hd__a21o_1 _07469_ (.A1(net1023),
    .A2(net343),
    .B1(_04075_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01867_));
 sky130_fd_sc_hd__mux2_1 _07470_ (.A0(\top.dut.bit_buf[5] ),
    .A1(net43),
    .S(net713),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04076_));
 sky130_fd_sc_hd__mux2_1 _07471_ (.A0(_04072_),
    .A1(_04076_),
    .S(_04049_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04077_));
 sky130_fd_sc_hd__mux2_1 _07472_ (.A0(_04055_),
    .A1(_04077_),
    .S(_04048_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04078_));
 sky130_fd_sc_hd__or2_1 _07473_ (.A(\top.dut.bits_in_buf_next[1] ),
    .B(_04052_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04079_));
 sky130_fd_sc_hd__o211a_1 _07474_ (.A1(net342),
    .A2(_04064_),
    .B1(_04079_),
    .C1(_04060_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04080_));
 sky130_fd_sc_hd__a221o_1 _07475_ (.A1(net1325),
    .A2(net344),
    .B1(_04045_),
    .B2(_04078_),
    .C1(_04080_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01866_));
 sky130_fd_sc_hd__mux2_1 _07476_ (.A0(\top.dut.bit_buf[4] ),
    .A1(net42),
    .S(net713),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04081_));
 sky130_fd_sc_hd__mux2_1 _07477_ (.A0(_04076_),
    .A1(_04081_),
    .S(net393),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04082_));
 sky130_fd_sc_hd__mux2_1 _07478_ (.A0(_04073_),
    .A1(_04082_),
    .S(net342),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04083_));
 sky130_fd_sc_hd__or2_1 _07479_ (.A(_04048_),
    .B(_04069_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04084_));
 sky130_fd_sc_hd__o211a_1 _07480_ (.A1(\top.dut.bits_in_buf_next[1] ),
    .A2(_04071_),
    .B1(_04084_),
    .C1(_04060_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04085_));
 sky130_fd_sc_hd__a221o_1 _07481_ (.A1(net1338),
    .A2(net344),
    .B1(_04045_),
    .B2(_04083_),
    .C1(_04085_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01865_));
 sky130_fd_sc_hd__mux2_1 _07482_ (.A0(\top.dut.bit_buf[3] ),
    .A1(net41),
    .S(net714),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04086_));
 sky130_fd_sc_hd__mux2_1 _07483_ (.A0(_04081_),
    .A1(_04086_),
    .S(net393),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04087_));
 sky130_fd_sc_hd__mux2_1 _07484_ (.A0(_04077_),
    .A1(_04087_),
    .S(net342),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04088_));
 sky130_fd_sc_hd__a22o_1 _07485_ (.A1(\top.dut.out[3] ),
    .A2(net344),
    .B1(_04056_),
    .B2(_04060_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04089_));
 sky130_fd_sc_hd__a21o_1 _07486_ (.A1(_04045_),
    .A2(_04088_),
    .B1(_04089_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01864_));
 sky130_fd_sc_hd__mux2_1 _07487_ (.A0(\top.dut.bit_buf[2] ),
    .A1(net40),
    .S(net713),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04090_));
 sky130_fd_sc_hd__mux2_1 _07488_ (.A0(_04086_),
    .A1(_04090_),
    .S(net393),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04091_));
 sky130_fd_sc_hd__mux2_1 _07489_ (.A0(_04082_),
    .A1(_04091_),
    .S(net342),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04092_));
 sky130_fd_sc_hd__a22o_1 _07490_ (.A1(\top.dut.out[2] ),
    .A2(net344),
    .B1(_04060_),
    .B2(_04074_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04093_));
 sky130_fd_sc_hd__a21o_1 _07491_ (.A1(_04045_),
    .A2(_04092_),
    .B1(_04093_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01863_));
 sky130_fd_sc_hd__mux2_1 _07492_ (.A0(\top.dut.bit_buf[1] ),
    .A1(net39),
    .S(net714),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04094_));
 sky130_fd_sc_hd__nor2_1 _07493_ (.A(\top.dut.bits_in_buf[1] ),
    .B(\top.dut.bits_in_buf_next[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04095_));
 sky130_fd_sc_hd__a32o_1 _07494_ (.A1(net342),
    .A2(\top.dut.bits_in_buf_next[0] ),
    .A3(_04090_),
    .B1(_04094_),
    .B2(_04095_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04096_));
 sky130_fd_sc_hd__a211o_1 _07495_ (.A1(\top.dut.bits_in_buf_next[1] ),
    .A2(_04087_),
    .B1(_04096_),
    .C1(_04046_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04097_));
 sky130_fd_sc_hd__o221a_1 _07496_ (.A1(net1620),
    .A2(\top.dut.out_valid_next ),
    .B1(_04061_),
    .B2(_04078_),
    .C1(_04097_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01862_));
 sky130_fd_sc_hd__mux2_1 _07497_ (.A0(\top.dut.bit_buf[0] ),
    .A1(net38),
    .S(net714),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04098_));
 sky130_fd_sc_hd__a221o_1 _07498_ (.A1(\top.dut.bits_in_buf_next[1] ),
    .A2(_04091_),
    .B1(_04095_),
    .B2(_04098_),
    .C1(_04046_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04099_));
 sky130_fd_sc_hd__a31o_1 _07499_ (.A1(net342),
    .A2(\top.dut.bits_in_buf_next[0] ),
    .A3(_04094_),
    .B1(_04099_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04100_));
 sky130_fd_sc_hd__o221a_1 _07500_ (.A1(net1628),
    .A2(\top.dut.out_valid_next ),
    .B1(_04061_),
    .B2(_04083_),
    .C1(_04100_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01861_));
 sky130_fd_sc_hd__a21o_1 _07501_ (.A1(_02980_),
    .A2(_02984_),
    .B1(_02982_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04101_));
 sky130_fd_sc_hd__a21oi_2 _07502_ (.A1(_02975_),
    .A2(_04101_),
    .B1(_02974_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04102_));
 sky130_fd_sc_hd__and2b_1 _07503_ (.A_N(_02990_),
    .B(_04102_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04103_));
 sky130_fd_sc_hd__nor2_2 _07504_ (.A(_02989_),
    .B(_04103_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04104_));
 sky130_fd_sc_hd__o31ai_2 _07505_ (.A1(_02979_),
    .A2(_02989_),
    .A3(_04103_),
    .B1(_02978_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04105_));
 sky130_fd_sc_hd__a21oi_1 _07506_ (.A1(_02988_),
    .A2(_04105_),
    .B1(_02986_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04106_));
 sky130_fd_sc_hd__xnor2_1 _07507_ (.A(_02972_),
    .B(_04106_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04107_));
 sky130_fd_sc_hd__xnor2_2 _07508_ (.A(_02988_),
    .B(_04105_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04108_));
 sky130_fd_sc_hd__xnor2_4 _07509_ (.A(_02979_),
    .B(_04104_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04109_));
 sky130_fd_sc_hd__xnor2_4 _07510_ (.A(_02991_),
    .B(_04102_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04110_));
 sky130_fd_sc_hd__xnor2_2 _07511_ (.A(_02975_),
    .B(_04101_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04111_));
 sky130_fd_sc_hd__xor2_1 _07512_ (.A(_02980_),
    .B(_02984_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04112_));
 sky130_fd_sc_hd__mux4_1 _07513_ (.A0(\top.cb_syn.char_path_n[110] ),
    .A1(\top.cb_syn.char_path_n[109] ),
    .A2(\top.cb_syn.char_path_n[112] ),
    .A3(\top.cb_syn.char_path_n[111] ),
    .S0(net396),
    .S1(net294),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04113_));
 sky130_fd_sc_hd__mux4_1 _07514_ (.A0(\top.cb_syn.char_path_n[106] ),
    .A1(\top.cb_syn.char_path_n[105] ),
    .A2(\top.cb_syn.char_path_n[108] ),
    .A3(\top.cb_syn.char_path_n[107] ),
    .S0(net395),
    .S1(net293),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04114_));
 sky130_fd_sc_hd__mux2_1 _07515_ (.A0(_04113_),
    .A1(_04114_),
    .S(net290),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04115_));
 sky130_fd_sc_hd__mux4_1 _07516_ (.A0(\top.cb_syn.char_path_n[102] ),
    .A1(\top.cb_syn.char_path_n[101] ),
    .A2(\top.cb_syn.char_path_n[104] ),
    .A3(\top.cb_syn.char_path_n[103] ),
    .S0(net395),
    .S1(net293),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04116_));
 sky130_fd_sc_hd__mux4_1 _07517_ (.A0(\top.cb_syn.char_path_n[98] ),
    .A1(\top.cb_syn.char_path_n[97] ),
    .A2(\top.cb_syn.char_path_n[100] ),
    .A3(\top.cb_syn.char_path_n[99] ),
    .S0(net395),
    .S1(net293),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04117_));
 sky130_fd_sc_hd__mux2_1 _07518_ (.A0(_04116_),
    .A1(_04117_),
    .S(net289),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04118_));
 sky130_fd_sc_hd__mux2_1 _07519_ (.A0(_04115_),
    .A1(_04118_),
    .S(_04110_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04119_));
 sky130_fd_sc_hd__mux4_1 _07520_ (.A0(\top.cb_syn.char_path_n[126] ),
    .A1(\top.cb_syn.char_path_n[125] ),
    .A2(\top.cb_syn.curr_path[127] ),
    .A3(\top.cb_syn.char_path_n[127] ),
    .S0(net394),
    .S1(net292),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04120_));
 sky130_fd_sc_hd__mux4_1 _07521_ (.A0(\top.cb_syn.char_path_n[122] ),
    .A1(\top.cb_syn.char_path_n[121] ),
    .A2(\top.cb_syn.char_path_n[124] ),
    .A3(\top.cb_syn.char_path_n[123] ),
    .S0(net394),
    .S1(net292),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04121_));
 sky130_fd_sc_hd__mux2_1 _07522_ (.A0(_04120_),
    .A1(_04121_),
    .S(net289),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04122_));
 sky130_fd_sc_hd__mux4_1 _07523_ (.A0(\top.cb_syn.char_path_n[118] ),
    .A1(\top.cb_syn.char_path_n[117] ),
    .A2(\top.cb_syn.char_path_n[120] ),
    .A3(\top.cb_syn.char_path_n[119] ),
    .S0(net394),
    .S1(net295),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04123_));
 sky130_fd_sc_hd__mux4_1 _07524_ (.A0(\top.cb_syn.char_path_n[114] ),
    .A1(\top.cb_syn.char_path_n[113] ),
    .A2(\top.cb_syn.char_path_n[116] ),
    .A3(\top.cb_syn.char_path_n[115] ),
    .S0(net396),
    .S1(net294),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04124_));
 sky130_fd_sc_hd__mux2_1 _07525_ (.A0(_04123_),
    .A1(_04124_),
    .S(net289),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04125_));
 sky130_fd_sc_hd__mux2_1 _07526_ (.A0(_04122_),
    .A1(_04125_),
    .S(_04110_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04126_));
 sky130_fd_sc_hd__mux2_1 _07527_ (.A0(_04119_),
    .A1(_04126_),
    .S(_04109_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04127_));
 sky130_fd_sc_hd__mux4_1 _07528_ (.A0(\top.cb_syn.char_path_n[78] ),
    .A1(\top.cb_syn.char_path_n[77] ),
    .A2(\top.cb_syn.char_path_n[80] ),
    .A3(\top.cb_syn.char_path_n[79] ),
    .S0(net397),
    .S1(net294),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04128_));
 sky130_fd_sc_hd__mux4_1 _07529_ (.A0(\top.cb_syn.char_path_n[74] ),
    .A1(\top.cb_syn.char_path_n[73] ),
    .A2(\top.cb_syn.char_path_n[76] ),
    .A3(\top.cb_syn.char_path_n[75] ),
    .S0(net397),
    .S1(net295),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04129_));
 sky130_fd_sc_hd__mux2_1 _07530_ (.A0(_04128_),
    .A1(_04129_),
    .S(net290),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04130_));
 sky130_fd_sc_hd__mux4_1 _07531_ (.A0(\top.cb_syn.char_path_n[70] ),
    .A1(\top.cb_syn.char_path_n[69] ),
    .A2(\top.cb_syn.char_path_n[72] ),
    .A3(\top.cb_syn.char_path_n[71] ),
    .S0(net395),
    .S1(net293),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04131_));
 sky130_fd_sc_hd__mux4_1 _07532_ (.A0(\top.cb_syn.char_path_n[66] ),
    .A1(\top.cb_syn.char_path_n[65] ),
    .A2(\top.cb_syn.char_path_n[68] ),
    .A3(\top.cb_syn.char_path_n[67] ),
    .S0(net395),
    .S1(net293),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04132_));
 sky130_fd_sc_hd__mux2_1 _07533_ (.A0(_04131_),
    .A1(_04132_),
    .S(net289),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04133_));
 sky130_fd_sc_hd__mux2_1 _07534_ (.A0(_04130_),
    .A1(_04133_),
    .S(_04110_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04134_));
 sky130_fd_sc_hd__mux4_1 _07535_ (.A0(\top.cb_syn.char_path_n[94] ),
    .A1(\top.cb_syn.char_path_n[93] ),
    .A2(\top.cb_syn.char_path_n[96] ),
    .A3(\top.cb_syn.char_path_n[95] ),
    .S0(net394),
    .S1(net292),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04135_));
 sky130_fd_sc_hd__mux4_1 _07536_ (.A0(\top.cb_syn.char_path_n[90] ),
    .A1(\top.cb_syn.char_path_n[89] ),
    .A2(\top.cb_syn.char_path_n[92] ),
    .A3(\top.cb_syn.char_path_n[91] ),
    .S0(net394),
    .S1(net292),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04136_));
 sky130_fd_sc_hd__mux2_1 _07537_ (.A0(_04135_),
    .A1(_04136_),
    .S(net289),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04137_));
 sky130_fd_sc_hd__mux4_1 _07538_ (.A0(\top.cb_syn.char_path_n[86] ),
    .A1(\top.cb_syn.char_path_n[85] ),
    .A2(\top.cb_syn.char_path_n[88] ),
    .A3(\top.cb_syn.char_path_n[87] ),
    .S0(net396),
    .S1(net294),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04138_));
 sky130_fd_sc_hd__mux4_1 _07539_ (.A0(\top.cb_syn.char_path_n[82] ),
    .A1(\top.cb_syn.char_path_n[81] ),
    .A2(\top.cb_syn.char_path_n[84] ),
    .A3(\top.cb_syn.char_path_n[83] ),
    .S0(net396),
    .S1(net294),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04139_));
 sky130_fd_sc_hd__mux2_1 _07540_ (.A0(_04138_),
    .A1(_04139_),
    .S(net289),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04140_));
 sky130_fd_sc_hd__mux2_1 _07541_ (.A0(_04137_),
    .A1(_04140_),
    .S(_04110_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04141_));
 sky130_fd_sc_hd__mux2_1 _07542_ (.A0(_04134_),
    .A1(_04141_),
    .S(_04109_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04142_));
 sky130_fd_sc_hd__mux2_1 _07543_ (.A0(_04127_),
    .A1(_04142_),
    .S(_04108_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04143_));
 sky130_fd_sc_hd__mux4_1 _07544_ (.A0(\top.cb_syn.char_path_n[14] ),
    .A1(\top.cb_syn.char_path_n[13] ),
    .A2(\top.cb_syn.char_path_n[16] ),
    .A3(\top.cb_syn.char_path_n[15] ),
    .S0(net395),
    .S1(net293),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04144_));
 sky130_fd_sc_hd__mux4_1 _07545_ (.A0(\top.cb_syn.char_path_n[10] ),
    .A1(\top.cb_syn.char_path_n[9] ),
    .A2(\top.cb_syn.char_path_n[12] ),
    .A3(\top.cb_syn.char_path_n[11] ),
    .S0(net396),
    .S1(net294),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04145_));
 sky130_fd_sc_hd__mux2_1 _07546_ (.A0(_04144_),
    .A1(_04145_),
    .S(net290),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04146_));
 sky130_fd_sc_hd__mux4_1 _07547_ (.A0(\top.cb_syn.char_path_n[6] ),
    .A1(\top.cb_syn.char_path_n[5] ),
    .A2(\top.cb_syn.char_path_n[8] ),
    .A3(\top.cb_syn.char_path_n[7] ),
    .S0(net396),
    .S1(net294),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04147_));
 sky130_fd_sc_hd__mux4_1 _07548_ (.A0(\top.cb_syn.char_path_n[2] ),
    .A1(\top.cb_syn.char_path_n[1] ),
    .A2(\top.cb_syn.char_path_n[4] ),
    .A3(\top.cb_syn.char_path_n[3] ),
    .S0(net396),
    .S1(net294),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04148_));
 sky130_fd_sc_hd__mux2_1 _07549_ (.A0(_04147_),
    .A1(_04148_),
    .S(net290),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04149_));
 sky130_fd_sc_hd__mux2_1 _07550_ (.A0(_04146_),
    .A1(_04149_),
    .S(_04110_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04150_));
 sky130_fd_sc_hd__mux4_1 _07551_ (.A0(\top.cb_syn.char_path_n[30] ),
    .A1(\top.cb_syn.char_path_n[29] ),
    .A2(\top.cb_syn.char_path_n[32] ),
    .A3(\top.cb_syn.char_path_n[31] ),
    .S0(net397),
    .S1(net292),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04151_));
 sky130_fd_sc_hd__mux4_1 _07552_ (.A0(\top.cb_syn.char_path_n[26] ),
    .A1(\top.cb_syn.char_path_n[25] ),
    .A2(\top.cb_syn.char_path_n[28] ),
    .A3(\top.cb_syn.char_path_n[27] ),
    .S0(net397),
    .S1(net292),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04152_));
 sky130_fd_sc_hd__mux2_1 _07553_ (.A0(_04151_),
    .A1(_04152_),
    .S(net289),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04153_));
 sky130_fd_sc_hd__mux4_1 _07554_ (.A0(\top.cb_syn.char_path_n[22] ),
    .A1(\top.cb_syn.char_path_n[21] ),
    .A2(\top.cb_syn.char_path_n[24] ),
    .A3(\top.cb_syn.char_path_n[23] ),
    .S0(net394),
    .S1(net292),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04154_));
 sky130_fd_sc_hd__mux4_1 _07555_ (.A0(\top.cb_syn.char_path_n[18] ),
    .A1(\top.cb_syn.char_path_n[17] ),
    .A2(\top.cb_syn.char_path_n[20] ),
    .A3(\top.cb_syn.char_path_n[19] ),
    .S0(net396),
    .S1(net294),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04155_));
 sky130_fd_sc_hd__mux2_1 _07556_ (.A0(_04154_),
    .A1(_04155_),
    .S(net289),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04156_));
 sky130_fd_sc_hd__mux2_1 _07557_ (.A0(_04153_),
    .A1(_04156_),
    .S(_04110_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04157_));
 sky130_fd_sc_hd__mux2_1 _07558_ (.A0(_04150_),
    .A1(_04157_),
    .S(_04109_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04158_));
 sky130_fd_sc_hd__mux4_1 _07559_ (.A0(\top.cb_syn.char_path_n[46] ),
    .A1(\top.cb_syn.char_path_n[45] ),
    .A2(\top.cb_syn.char_path_n[48] ),
    .A3(\top.cb_syn.char_path_n[47] ),
    .S0(net395),
    .S1(net293),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04159_));
 sky130_fd_sc_hd__mux4_1 _07560_ (.A0(\top.cb_syn.char_path_n[42] ),
    .A1(\top.cb_syn.char_path_n[41] ),
    .A2(\top.cb_syn.char_path_n[44] ),
    .A3(\top.cb_syn.char_path_n[43] ),
    .S0(net395),
    .S1(net293),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04160_));
 sky130_fd_sc_hd__mux2_1 _07561_ (.A0(_04159_),
    .A1(_04160_),
    .S(net290),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04161_));
 sky130_fd_sc_hd__mux4_1 _07562_ (.A0(\top.cb_syn.char_path_n[38] ),
    .A1(\top.cb_syn.char_path_n[37] ),
    .A2(\top.cb_syn.char_path_n[40] ),
    .A3(\top.cb_syn.char_path_n[39] ),
    .S0(net395),
    .S1(net293),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04162_));
 sky130_fd_sc_hd__mux4_1 _07563_ (.A0(\top.cb_syn.char_path_n[34] ),
    .A1(\top.cb_syn.char_path_n[33] ),
    .A2(\top.cb_syn.char_path_n[36] ),
    .A3(\top.cb_syn.char_path_n[35] ),
    .S0(net395),
    .S1(net293),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04163_));
 sky130_fd_sc_hd__mux2_1 _07564_ (.A0(_04162_),
    .A1(_04163_),
    .S(net290),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04164_));
 sky130_fd_sc_hd__mux2_1 _07565_ (.A0(_04161_),
    .A1(_04164_),
    .S(_04110_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04165_));
 sky130_fd_sc_hd__mux4_1 _07566_ (.A0(\top.cb_syn.char_path_n[62] ),
    .A1(\top.cb_syn.char_path_n[61] ),
    .A2(\top.cb_syn.char_path_n[64] ),
    .A3(\top.cb_syn.char_path_n[63] ),
    .S0(net394),
    .S1(net292),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04166_));
 sky130_fd_sc_hd__mux4_1 _07567_ (.A0(\top.cb_syn.char_path_n[58] ),
    .A1(\top.cb_syn.char_path_n[57] ),
    .A2(\top.cb_syn.char_path_n[60] ),
    .A3(\top.cb_syn.char_path_n[59] ),
    .S0(net394),
    .S1(net292),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04167_));
 sky130_fd_sc_hd__mux2_1 _07568_ (.A0(_04166_),
    .A1(_04167_),
    .S(net289),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04168_));
 sky130_fd_sc_hd__mux4_1 _07569_ (.A0(\top.cb_syn.char_path_n[54] ),
    .A1(\top.cb_syn.char_path_n[53] ),
    .A2(\top.cb_syn.char_path_n[56] ),
    .A3(\top.cb_syn.char_path_n[55] ),
    .S0(net394),
    .S1(net295),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04169_));
 sky130_fd_sc_hd__mux4_1 _07570_ (.A0(\top.cb_syn.char_path_n[50] ),
    .A1(\top.cb_syn.char_path_n[49] ),
    .A2(\top.cb_syn.char_path_n[52] ),
    .A3(\top.cb_syn.char_path_n[51] ),
    .S0(net396),
    .S1(net292),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04170_));
 sky130_fd_sc_hd__mux2_1 _07571_ (.A0(_04169_),
    .A1(_04170_),
    .S(net289),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04171_));
 sky130_fd_sc_hd__mux2_1 _07572_ (.A0(_04168_),
    .A1(_04171_),
    .S(_04110_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04172_));
 sky130_fd_sc_hd__mux2_1 _07573_ (.A0(_04165_),
    .A1(_04172_),
    .S(_04109_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04173_));
 sky130_fd_sc_hd__mux2_1 _07574_ (.A0(_04173_),
    .A1(_04158_),
    .S(_04108_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04174_));
 sky130_fd_sc_hd__mux2_1 _07575_ (.A0(_04143_),
    .A1(_04174_),
    .S(_04107_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04175_));
 sky130_fd_sc_hd__or2_4 _07576_ (.A(_02551_),
    .B(_04175_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04176_));
 sky130_fd_sc_hd__mux2_1 _07577_ (.A0(\top.cb_syn.h_element[61] ),
    .A1(\top.cb_syn.h_element[52] ),
    .S(_04176_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04177_));
 sky130_fd_sc_hd__or2_2 _07578_ (.A(net519),
    .B(net524),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04178_));
 sky130_fd_sc_hd__or2_2 _07579_ (.A(net516),
    .B(net521),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04179_));
 sky130_fd_sc_hd__nor2_2 _07580_ (.A(_04178_),
    .B(_04179_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04180_));
 sky130_fd_sc_hd__or2_2 _07581_ (.A(_04178_),
    .B(_04179_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04181_));
 sky130_fd_sc_hd__a221o_1 _07582_ (.A1(net517),
    .A2(\top.cb_syn.h_element[52] ),
    .B1(net525),
    .B2(\top.cb_syn.h_element[61] ),
    .C1(_04180_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04182_));
 sky130_fd_sc_hd__or3_1 _07583_ (.A(\top.cb_syn.max_index[3] ),
    .B(\top.cb_syn.max_index[2] ),
    .C(\top.cb_syn.max_index[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04183_));
 sky130_fd_sc_hd__or2_1 _07584_ (.A(\top.cb_syn.max_index[4] ),
    .B(_04183_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04184_));
 sky130_fd_sc_hd__or3_1 _07585_ (.A(\top.cb_syn.max_index[6] ),
    .B(\top.cb_syn.max_index[5] ),
    .C(_04184_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04185_));
 sky130_fd_sc_hd__xnor2_1 _07586_ (.A(\top.cb_syn.max_index[7] ),
    .B(_04185_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04186_));
 sky130_fd_sc_hd__a22o_1 _07587_ (.A1(net521),
    .A2(_04177_),
    .B1(_04186_),
    .B2(net516),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04187_));
 sky130_fd_sc_hd__o21a_1 _07588_ (.A1(_02972_),
    .A2(_04106_),
    .B1(_02971_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04188_));
 sky130_fd_sc_hd__nor2_1 _07589_ (.A(_02993_),
    .B(_04188_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04189_));
 sky130_fd_sc_hd__or2_2 _07590_ (.A(\top.cb_syn.pulse_first ),
    .B(_02891_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04190_));
 sky130_fd_sc_hd__inv_2 _07591_ (.A(_04190_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04191_));
 sky130_fd_sc_hd__nor2_1 _07592_ (.A(\top.cb_syn.h_element[54] ),
    .B(_04190_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04192_));
 sky130_fd_sc_hd__and4_1 _07593_ (.A(net550),
    .B(_04175_),
    .C(_04189_),
    .D(_04192_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04193_));
 sky130_fd_sc_hd__a21oi_1 _07594_ (.A1(net550),
    .A2(_04189_),
    .B1(_04190_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04194_));
 sky130_fd_sc_hd__nand2_1 _07595_ (.A(net519),
    .B(_02884_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04195_));
 sky130_fd_sc_hd__o21a_1 _07596_ (.A1(net412),
    .A2(_02884_),
    .B1(_02886_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04196_));
 sky130_fd_sc_hd__and2_1 _07597_ (.A(net412),
    .B(_02896_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04197_));
 sky130_fd_sc_hd__or3_1 _07598_ (.A(\top.cb_syn.cb_length[4] ),
    .B(\top.cb_syn.cb_length[3] ),
    .C(\top.cb_syn.cb_length[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04198_));
 sky130_fd_sc_hd__or3_1 _07599_ (.A(\top.cb_syn.cb_length[6] ),
    .B(\top.cb_syn.cb_length[5] ),
    .C(_04198_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04199_));
 sky130_fd_sc_hd__or3_1 _07600_ (.A(\top.cb_syn.cb_length[2] ),
    .B(\top.cb_syn.cb_length[1] ),
    .C(\top.cb_syn.cb_length[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04200_));
 sky130_fd_sc_hd__or3_2 _07601_ (.A(\top.cb_syn.cb_length[1] ),
    .B(\top.cb_syn.cb_length[0] ),
    .C(_04199_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04201_));
 sky130_fd_sc_hd__nor2_1 _07602_ (.A(_02543_),
    .B(_04201_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04202_));
 sky130_fd_sc_hd__or3b_1 _07603_ (.A(net489),
    .B(_02895_),
    .C_N(net524),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04203_));
 sky130_fd_sc_hd__and3_1 _07604_ (.A(\top.cb_syn.pulse_first ),
    .B(net521),
    .C(_02889_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04204_));
 sky130_fd_sc_hd__a221o_1 _07605_ (.A1(_02525_),
    .A2(\top.cb_syn.curr_state[0] ),
    .B1(_04178_),
    .B2(net488),
    .C1(_04204_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04205_));
 sky130_fd_sc_hd__or2_1 _07606_ (.A(net488),
    .B(net423),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04206_));
 sky130_fd_sc_hd__a21o_1 _07607_ (.A1(net522),
    .A2(_02890_),
    .B1(net423),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04207_));
 sky130_fd_sc_hd__inv_2 _07608_ (.A(_04207_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04208_));
 sky130_fd_sc_hd__nor2_1 _07609_ (.A(\top.cb_syn.curr_state[0] ),
    .B(_04181_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04209_));
 sky130_fd_sc_hd__or4b_1 _07610_ (.A(_04205_),
    .B(_04207_),
    .C(_04209_),
    .D_N(_04203_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04210_));
 sky130_fd_sc_hd__or4_1 _07611_ (.A(_04196_),
    .B(_04197_),
    .C(_04202_),
    .D(_04210_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04211_));
 sky130_fd_sc_hd__nor3_4 _07612_ (.A(_04193_),
    .B(_04194_),
    .C(_04211_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04212_));
 sky130_fd_sc_hd__o22a_1 _07613_ (.A1(\top.cb_syn.max_index[7] ),
    .A2(_04181_),
    .B1(_04182_),
    .B2(_04187_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04213_));
 sky130_fd_sc_hd__mux2_1 _07614_ (.A0(net1499),
    .A1(_04213_),
    .S(_04212_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01860_));
 sky130_fd_sc_hd__mux2_1 _07615_ (.A0(\top.cb_syn.h_element[60] ),
    .A1(\top.cb_syn.h_element[51] ),
    .S(_04176_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04214_));
 sky130_fd_sc_hd__a221o_1 _07616_ (.A1(net518),
    .A2(\top.cb_syn.h_element[51] ),
    .B1(net525),
    .B2(\top.cb_syn.h_element[60] ),
    .C1(_04180_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04215_));
 sky130_fd_sc_hd__o21ai_1 _07617_ (.A1(\top.cb_syn.max_index[5] ),
    .A2(_04184_),
    .B1(\top.cb_syn.max_index[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04216_));
 sky130_fd_sc_hd__nand2_1 _07618_ (.A(_04185_),
    .B(_04216_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04217_));
 sky130_fd_sc_hd__a22o_1 _07619_ (.A1(net521),
    .A2(_04214_),
    .B1(_04217_),
    .B2(net516),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04218_));
 sky130_fd_sc_hd__o22a_1 _07620_ (.A1(\top.cb_syn.max_index[6] ),
    .A2(_04181_),
    .B1(_04215_),
    .B2(_04218_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04219_));
 sky130_fd_sc_hd__mux2_1 _07621_ (.A0(net1417),
    .A1(_04219_),
    .S(_04212_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01859_));
 sky130_fd_sc_hd__mux2_1 _07622_ (.A0(\top.cb_syn.h_element[59] ),
    .A1(\top.cb_syn.h_element[50] ),
    .S(_04176_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04220_));
 sky130_fd_sc_hd__a221o_1 _07623_ (.A1(net517),
    .A2(\top.cb_syn.h_element[50] ),
    .B1(net525),
    .B2(\top.cb_syn.h_element[59] ),
    .C1(_04180_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04221_));
 sky130_fd_sc_hd__xnor2_1 _07624_ (.A(\top.cb_syn.max_index[5] ),
    .B(_04184_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04222_));
 sky130_fd_sc_hd__a22o_1 _07625_ (.A1(net521),
    .A2(_04220_),
    .B1(_04222_),
    .B2(net516),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04223_));
 sky130_fd_sc_hd__o22a_1 _07626_ (.A1(\top.cb_syn.max_index[5] ),
    .A2(_04181_),
    .B1(_04221_),
    .B2(_04223_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04224_));
 sky130_fd_sc_hd__mux2_1 _07627_ (.A0(net1550),
    .A1(_04224_),
    .S(_04212_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01858_));
 sky130_fd_sc_hd__mux2_1 _07628_ (.A0(\top.cb_syn.h_element[58] ),
    .A1(\top.cb_syn.h_element[49] ),
    .S(_04176_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04225_));
 sky130_fd_sc_hd__a221o_1 _07629_ (.A1(net517),
    .A2(\top.cb_syn.h_element[49] ),
    .B1(net525),
    .B2(\top.cb_syn.h_element[58] ),
    .C1(_04180_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04226_));
 sky130_fd_sc_hd__nand2_1 _07630_ (.A(\top.cb_syn.max_index[4] ),
    .B(_04183_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04227_));
 sky130_fd_sc_hd__nand2_1 _07631_ (.A(_04184_),
    .B(_04227_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04228_));
 sky130_fd_sc_hd__a22o_1 _07632_ (.A1(net521),
    .A2(_04225_),
    .B1(_04228_),
    .B2(net516),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04229_));
 sky130_fd_sc_hd__o22a_1 _07633_ (.A1(\top.cb_syn.max_index[4] ),
    .A2(_04181_),
    .B1(_04226_),
    .B2(_04229_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04230_));
 sky130_fd_sc_hd__mux2_1 _07634_ (.A0(net1500),
    .A1(_04230_),
    .S(_04212_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01857_));
 sky130_fd_sc_hd__mux2_1 _07635_ (.A0(\top.cb_syn.h_element[57] ),
    .A1(\top.cb_syn.h_element[48] ),
    .S(_04176_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04231_));
 sky130_fd_sc_hd__a221o_1 _07636_ (.A1(net518),
    .A2(\top.cb_syn.h_element[48] ),
    .B1(net525),
    .B2(\top.cb_syn.h_element[57] ),
    .C1(_04180_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04232_));
 sky130_fd_sc_hd__o21ai_1 _07637_ (.A1(\top.cb_syn.max_index[2] ),
    .A2(\top.cb_syn.max_index[1] ),
    .B1(\top.cb_syn.max_index[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04233_));
 sky130_fd_sc_hd__nand2_1 _07638_ (.A(_04183_),
    .B(_04233_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04234_));
 sky130_fd_sc_hd__a22o_1 _07639_ (.A1(net521),
    .A2(_04231_),
    .B1(_04234_),
    .B2(net516),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04235_));
 sky130_fd_sc_hd__o22a_1 _07640_ (.A1(\top.cb_syn.max_index[3] ),
    .A2(_04181_),
    .B1(_04232_),
    .B2(_04235_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04236_));
 sky130_fd_sc_hd__mux2_1 _07641_ (.A0(net1455),
    .A1(_04236_),
    .S(_04212_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01856_));
 sky130_fd_sc_hd__mux2_1 _07642_ (.A0(\top.cb_syn.h_element[56] ),
    .A1(\top.cb_syn.h_element[47] ),
    .S(_04176_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04237_));
 sky130_fd_sc_hd__a221o_1 _07643_ (.A1(net518),
    .A2(\top.cb_syn.h_element[47] ),
    .B1(net525),
    .B2(\top.cb_syn.h_element[56] ),
    .C1(_04180_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04238_));
 sky130_fd_sc_hd__xor2_1 _07644_ (.A(\top.cb_syn.max_index[2] ),
    .B(\top.cb_syn.max_index[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04239_));
 sky130_fd_sc_hd__inv_2 _07645_ (.A(_04239_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04240_));
 sky130_fd_sc_hd__a22o_1 _07646_ (.A1(net521),
    .A2(_04237_),
    .B1(_04240_),
    .B2(net516),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04241_));
 sky130_fd_sc_hd__o22a_1 _07647_ (.A1(\top.cb_syn.max_index[2] ),
    .A2(_04181_),
    .B1(_04238_),
    .B2(_04241_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04242_));
 sky130_fd_sc_hd__mux2_1 _07648_ (.A0(net1070),
    .A1(_04242_),
    .S(_04212_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01855_));
 sky130_fd_sc_hd__mux2_1 _07649_ (.A0(\top.cb_syn.h_element[55] ),
    .A1(\top.cb_syn.h_element[46] ),
    .S(_04176_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04243_));
 sky130_fd_sc_hd__a2bb2o_1 _07650_ (.A1_N(_02543_),
    .A2_N(\top.cb_syn.max_index[1] ),
    .B1(\top.cb_syn.h_element[46] ),
    .B2(net517),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04244_));
 sky130_fd_sc_hd__a221o_1 _07651_ (.A1(\top.cb_syn.h_element[55] ),
    .A2(net525),
    .B1(_04180_),
    .B2(\top.cb_syn.max_index[1] ),
    .C1(_04244_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04245_));
 sky130_fd_sc_hd__a21o_1 _07652_ (.A1(net521),
    .A2(_04243_),
    .B1(_04245_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04246_));
 sky130_fd_sc_hd__mux2_1 _07653_ (.A0(net1556),
    .A1(_04246_),
    .S(_04212_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01854_));
 sky130_fd_sc_hd__or2_1 _07654_ (.A(_02831_),
    .B(_02835_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04247_));
 sky130_fd_sc_hd__nand3_4 _07655_ (.A(_02837_),
    .B(_02853_),
    .C(_04247_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04248_));
 sky130_fd_sc_hd__and4_2 _07656_ (.A(\top.findLeastValue.least2[8] ),
    .B(\top.findLeastValue.least1[8] ),
    .C(_02837_),
    .D(_04247_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04249_));
 sky130_fd_sc_hd__a21o_1 _07657_ (.A1(net449),
    .A2(net282),
    .B1(net1000),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01853_));
 sky130_fd_sc_hd__or2_1 _07658_ (.A(\top.hTree.write_HT_fin ),
    .B(\top.hTree.closing ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04250_));
 sky130_fd_sc_hd__nand2_2 _07659_ (.A(_04248_),
    .B(net388),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04251_));
 sky130_fd_sc_hd__o22ai_1 _07660_ (.A1(\top.findLeastValue.least1[8] ),
    .A2(net390),
    .B1(net265),
    .B2(\top.hTree.tree_reg[63] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04252_));
 sky130_fd_sc_hd__nand2_1 _07661_ (.A(net471),
    .B(_04252_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04253_));
 sky130_fd_sc_hd__nor2_2 _07662_ (.A(\top.hTree.write_HT_fin ),
    .B(_02837_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04254_));
 sky130_fd_sc_hd__or2_4 _07663_ (.A(\top.hTree.write_HT_fin ),
    .B(_02837_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04255_));
 sky130_fd_sc_hd__nor2_2 _07664_ (.A(net433),
    .B(_04254_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04256_));
 sky130_fd_sc_hd__nand2_4 _07665_ (.A(net449),
    .B(_04255_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04257_));
 sky130_fd_sc_hd__or3_1 _07666_ (.A(\top.hTree.tree_reg[63] ),
    .B(net471),
    .C(net282),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04258_));
 sky130_fd_sc_hd__a32o_1 _07667_ (.A1(_04253_),
    .A2(net256),
    .A3(_04258_),
    .B1(net1371),
    .B2(net431),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01852_));
 sky130_fd_sc_hd__mux2_1 _07668_ (.A0(\top.findLeastValue.least1[7] ),
    .A1(\top.hTree.tree_reg[62] ),
    .S(_04248_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04259_));
 sky130_fd_sc_hd__mux2_1 _07669_ (.A0(\top.findLeastValue.least1[7] ),
    .A1(_04259_),
    .S(net389),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04260_));
 sky130_fd_sc_hd__mux2_1 _07670_ (.A0(_04259_),
    .A1(_04260_),
    .S(net474),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04261_));
 sky130_fd_sc_hd__o22a_1 _07671_ (.A1(net449),
    .A2(net1160),
    .B1(_04257_),
    .B2(_04261_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01851_));
 sky130_fd_sc_hd__mux2_1 _07672_ (.A0(\top.findLeastValue.least1[6] ),
    .A1(\top.hTree.tree_reg[61] ),
    .S(_04248_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04262_));
 sky130_fd_sc_hd__mux2_1 _07673_ (.A0(\top.findLeastValue.least1[6] ),
    .A1(_04262_),
    .S(net389),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04263_));
 sky130_fd_sc_hd__mux2_1 _07674_ (.A0(_04262_),
    .A1(_04263_),
    .S(net474),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04264_));
 sky130_fd_sc_hd__o22a_1 _07675_ (.A1(net449),
    .A2(net1039),
    .B1(_04257_),
    .B2(_04264_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01850_));
 sky130_fd_sc_hd__and3_1 _07676_ (.A(\top.hTree.tree_reg[60] ),
    .B(_04248_),
    .C(net387),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04265_));
 sky130_fd_sc_hd__mux2_1 _07677_ (.A0(\top.hTree.tree_reg[60] ),
    .A1(\top.findLeastValue.least1[5] ),
    .S(net280),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04266_));
 sky130_fd_sc_hd__a21oi_1 _07678_ (.A1(\top.findLeastValue.least1[5] ),
    .A2(net264),
    .B1(_04265_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04267_));
 sky130_fd_sc_hd__nand2_1 _07679_ (.A(net472),
    .B(_04267_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04268_));
 sky130_fd_sc_hd__or2_1 _07680_ (.A(net472),
    .B(_04266_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04269_));
 sky130_fd_sc_hd__a32o_1 _07681_ (.A1(net257),
    .A2(_04268_),
    .A3(_04269_),
    .B1(net1131),
    .B2(net433),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01849_));
 sky130_fd_sc_hd__and3_1 _07682_ (.A(\top.hTree.tree_reg[59] ),
    .B(_04248_),
    .C(net389),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04270_));
 sky130_fd_sc_hd__mux2_1 _07683_ (.A0(\top.hTree.tree_reg[59] ),
    .A1(\top.findLeastValue.least1[4] ),
    .S(net280),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04271_));
 sky130_fd_sc_hd__a21oi_1 _07684_ (.A1(\top.findLeastValue.least1[4] ),
    .A2(net264),
    .B1(_04270_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04272_));
 sky130_fd_sc_hd__nand2_1 _07685_ (.A(net474),
    .B(_04272_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04273_));
 sky130_fd_sc_hd__or2_1 _07686_ (.A(net474),
    .B(_04271_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04274_));
 sky130_fd_sc_hd__a32o_1 _07687_ (.A1(net257),
    .A2(_04273_),
    .A3(_04274_),
    .B1(net1195),
    .B2(net432),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01848_));
 sky130_fd_sc_hd__and3_1 _07688_ (.A(\top.hTree.tree_reg[58] ),
    .B(_04248_),
    .C(net389),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04275_));
 sky130_fd_sc_hd__mux2_1 _07689_ (.A0(\top.hTree.tree_reg[58] ),
    .A1(\top.findLeastValue.least1[3] ),
    .S(net280),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04276_));
 sky130_fd_sc_hd__a21oi_1 _07690_ (.A1(\top.findLeastValue.least1[3] ),
    .A2(net264),
    .B1(_04275_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04277_));
 sky130_fd_sc_hd__nand2_1 _07691_ (.A(net474),
    .B(_04277_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04278_));
 sky130_fd_sc_hd__or2_1 _07692_ (.A(net474),
    .B(_04276_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04279_));
 sky130_fd_sc_hd__a32o_1 _07693_ (.A1(net258),
    .A2(_04278_),
    .A3(_04279_),
    .B1(net1092),
    .B2(net432),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01847_));
 sky130_fd_sc_hd__and3_1 _07694_ (.A(\top.hTree.tree_reg[57] ),
    .B(_04248_),
    .C(net388),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04280_));
 sky130_fd_sc_hd__mux2_1 _07695_ (.A0(\top.hTree.tree_reg[57] ),
    .A1(\top.findLeastValue.least1[2] ),
    .S(net280),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04281_));
 sky130_fd_sc_hd__a21oi_1 _07696_ (.A1(\top.findLeastValue.least1[2] ),
    .A2(net264),
    .B1(_04280_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04282_));
 sky130_fd_sc_hd__nand2_1 _07697_ (.A(net473),
    .B(_04282_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04283_));
 sky130_fd_sc_hd__or2_1 _07698_ (.A(net473),
    .B(_04281_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04284_));
 sky130_fd_sc_hd__a32o_1 _07699_ (.A1(net257),
    .A2(_04283_),
    .A3(_04284_),
    .B1(net1073),
    .B2(net432),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01846_));
 sky130_fd_sc_hd__and3_1 _07700_ (.A(\top.hTree.tree_reg[56] ),
    .B(_04248_),
    .C(net388),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04285_));
 sky130_fd_sc_hd__mux2_1 _07701_ (.A0(\top.hTree.tree_reg[56] ),
    .A1(\top.findLeastValue.least1[1] ),
    .S(net281),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04286_));
 sky130_fd_sc_hd__a21oi_1 _07702_ (.A1(\top.findLeastValue.least1[1] ),
    .A2(net264),
    .B1(_04285_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04287_));
 sky130_fd_sc_hd__nand2_1 _07703_ (.A(net473),
    .B(_04287_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04288_));
 sky130_fd_sc_hd__or2_1 _07704_ (.A(net473),
    .B(_04286_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04289_));
 sky130_fd_sc_hd__a32o_1 _07705_ (.A1(net257),
    .A2(_04288_),
    .A3(_04289_),
    .B1(net1191),
    .B2(net432),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01845_));
 sky130_fd_sc_hd__and3_1 _07706_ (.A(\top.hTree.tree_reg[55] ),
    .B(_04248_),
    .C(net387),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04290_));
 sky130_fd_sc_hd__mux2_1 _07707_ (.A0(\top.hTree.tree_reg[55] ),
    .A1(\top.findLeastValue.least1[0] ),
    .S(net280),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04291_));
 sky130_fd_sc_hd__a21oi_1 _07708_ (.A1(\top.findLeastValue.least1[0] ),
    .A2(net264),
    .B1(_04290_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04292_));
 sky130_fd_sc_hd__nand2_1 _07709_ (.A(net475),
    .B(_04292_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04293_));
 sky130_fd_sc_hd__or2_1 _07710_ (.A(net475),
    .B(_04291_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04294_));
 sky130_fd_sc_hd__a32o_1 _07711_ (.A1(net258),
    .A2(_04293_),
    .A3(_04294_),
    .B1(net1175),
    .B2(net432),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01844_));
 sky130_fd_sc_hd__o221a_1 _07712_ (.A1(\top.findLeastValue.least2[8] ),
    .A2(net390),
    .B1(net265),
    .B2(\top.hTree.tree_reg[54] ),
    .C1(net470),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04295_));
 sky130_fd_sc_hd__o21a_1 _07713_ (.A1(\top.hTree.tree_reg[54] ),
    .A2(net282),
    .B1(net417),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04296_));
 sky130_fd_sc_hd__o32a_1 _07714_ (.A1(_04257_),
    .A2(_04295_),
    .A3(_04296_),
    .B1(net1619),
    .B2(net449),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01843_));
 sky130_fd_sc_hd__mux2_1 _07715_ (.A0(\top.findLeastValue.least2[7] ),
    .A1(\top.hTree.tree_reg[53] ),
    .S(_04248_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04297_));
 sky130_fd_sc_hd__mux2_1 _07716_ (.A0(\top.findLeastValue.least2[7] ),
    .A1(_04297_),
    .S(net389),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04298_));
 sky130_fd_sc_hd__mux2_1 _07717_ (.A0(_04297_),
    .A1(_04298_),
    .S(net474),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04299_));
 sky130_fd_sc_hd__o22a_1 _07718_ (.A1(net449),
    .A2(net1066),
    .B1(_04257_),
    .B2(_04299_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01842_));
 sky130_fd_sc_hd__mux2_1 _07719_ (.A0(\top.hTree.tree_reg[52] ),
    .A1(\top.findLeastValue.least2[6] ),
    .S(net280),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04300_));
 sky130_fd_sc_hd__nand2_1 _07720_ (.A(net387),
    .B(_04300_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04301_));
 sky130_fd_sc_hd__o21a_1 _07721_ (.A1(_02515_),
    .A2(net387),
    .B1(_04301_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04302_));
 sky130_fd_sc_hd__nand2_1 _07722_ (.A(net472),
    .B(_04302_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04303_));
 sky130_fd_sc_hd__or2_1 _07723_ (.A(net472),
    .B(_04300_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04304_));
 sky130_fd_sc_hd__a32o_1 _07724_ (.A1(net257),
    .A2(_04303_),
    .A3(_04304_),
    .B1(net1009),
    .B2(net432),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01841_));
 sky130_fd_sc_hd__mux2_1 _07725_ (.A0(\top.hTree.tree_reg[51] ),
    .A1(\top.findLeastValue.least2[5] ),
    .S(net280),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04305_));
 sky130_fd_sc_hd__nand2_1 _07726_ (.A(net387),
    .B(_04305_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04306_));
 sky130_fd_sc_hd__o21a_1 _07727_ (.A1(_02516_),
    .A2(net387),
    .B1(_04306_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04307_));
 sky130_fd_sc_hd__nand2_1 _07728_ (.A(net472),
    .B(_04307_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04308_));
 sky130_fd_sc_hd__or2_1 _07729_ (.A(net472),
    .B(_04305_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04309_));
 sky130_fd_sc_hd__a32o_1 _07730_ (.A1(net257),
    .A2(_04308_),
    .A3(_04309_),
    .B1(net985),
    .B2(net433),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01840_));
 sky130_fd_sc_hd__mux2_1 _07731_ (.A0(\top.hTree.tree_reg[50] ),
    .A1(\top.findLeastValue.least2[4] ),
    .S(net280),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04310_));
 sky130_fd_sc_hd__nand2_1 _07732_ (.A(net388),
    .B(_04310_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04311_));
 sky130_fd_sc_hd__o21a_1 _07733_ (.A1(_02517_),
    .A2(net388),
    .B1(_04311_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04312_));
 sky130_fd_sc_hd__nand2_1 _07734_ (.A(net473),
    .B(_04312_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04313_));
 sky130_fd_sc_hd__or2_1 _07735_ (.A(net473),
    .B(_04310_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04314_));
 sky130_fd_sc_hd__a32o_1 _07736_ (.A1(net257),
    .A2(_04313_),
    .A3(_04314_),
    .B1(net994),
    .B2(net432),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01839_));
 sky130_fd_sc_hd__mux2_1 _07737_ (.A0(\top.hTree.tree_reg[49] ),
    .A1(\top.findLeastValue.least2[3] ),
    .S(net280),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04315_));
 sky130_fd_sc_hd__nand2_1 _07738_ (.A(net389),
    .B(_04315_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04316_));
 sky130_fd_sc_hd__o21a_1 _07739_ (.A1(_02518_),
    .A2(net389),
    .B1(_04316_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04317_));
 sky130_fd_sc_hd__nand2_1 _07740_ (.A(net474),
    .B(_04317_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04318_));
 sky130_fd_sc_hd__or2_1 _07741_ (.A(net473),
    .B(_04315_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04319_));
 sky130_fd_sc_hd__a32o_1 _07742_ (.A1(net257),
    .A2(_04318_),
    .A3(_04319_),
    .B1(net1010),
    .B2(net432),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01838_));
 sky130_fd_sc_hd__mux2_1 _07743_ (.A0(\top.hTree.tree_reg[48] ),
    .A1(\top.findLeastValue.least2[2] ),
    .S(net280),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04320_));
 sky130_fd_sc_hd__nand2_1 _07744_ (.A(net387),
    .B(_04320_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04321_));
 sky130_fd_sc_hd__o21a_1 _07745_ (.A1(_02519_),
    .A2(net387),
    .B1(_04321_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04322_));
 sky130_fd_sc_hd__nand2_1 _07746_ (.A(net472),
    .B(_04322_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04323_));
 sky130_fd_sc_hd__or2_1 _07747_ (.A(net472),
    .B(_04320_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04324_));
 sky130_fd_sc_hd__a32o_1 _07748_ (.A1(net257),
    .A2(_04323_),
    .A3(_04324_),
    .B1(net997),
    .B2(net433),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01837_));
 sky130_fd_sc_hd__mux2_1 _07749_ (.A0(\top.hTree.tree_reg[47] ),
    .A1(\top.findLeastValue.least2[1] ),
    .S(net281),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04325_));
 sky130_fd_sc_hd__nand2_1 _07750_ (.A(net387),
    .B(_04325_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04326_));
 sky130_fd_sc_hd__o21a_1 _07751_ (.A1(_02520_),
    .A2(net387),
    .B1(_04326_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04327_));
 sky130_fd_sc_hd__nand2_1 _07752_ (.A(net472),
    .B(_04327_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04328_));
 sky130_fd_sc_hd__or2_1 _07753_ (.A(net472),
    .B(_04325_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04329_));
 sky130_fd_sc_hd__a32o_1 _07754_ (.A1(net257),
    .A2(_04328_),
    .A3(_04329_),
    .B1(net1011),
    .B2(net433),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01836_));
 sky130_fd_sc_hd__mux2_1 _07755_ (.A0(\top.hTree.tree_reg[46] ),
    .A1(\top.findLeastValue.least2[0] ),
    .S(net281),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04330_));
 sky130_fd_sc_hd__mux2_1 _07756_ (.A0(\top.hTree.tree_reg[46] ),
    .A1(\top.findLeastValue.least2[0] ),
    .S(net264),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04331_));
 sky130_fd_sc_hd__mux2_1 _07757_ (.A0(_04330_),
    .A1(_04331_),
    .S(net475),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04332_));
 sky130_fd_sc_hd__a22o_1 _07758_ (.A1(net433),
    .A2(net1510),
    .B1(net258),
    .B2(_04332_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01835_));
 sky130_fd_sc_hd__mux2_1 _07759_ (.A0(\top.hTree.tree_reg[45] ),
    .A1(\top.findLeastValue.sum[45] ),
    .S(net286),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04333_));
 sky130_fd_sc_hd__mux2_1 _07760_ (.A0(\top.hTree.tree_reg[45] ),
    .A1(\top.findLeastValue.sum[45] ),
    .S(net267),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04334_));
 sky130_fd_sc_hd__or2_1 _07761_ (.A(net478),
    .B(_04333_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04335_));
 sky130_fd_sc_hd__o211a_1 _07762_ (.A1(net421),
    .A2(_04334_),
    .B1(_04335_),
    .C1(net263),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04336_));
 sky130_fd_sc_hd__nor2_1 _07763_ (.A(net431),
    .B(_04255_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04337_));
 sky130_fd_sc_hd__a221o_1 _07764_ (.A1(net438),
    .A2(net1582),
    .B1(net252),
    .B2(\top.findLeastValue.sum[45] ),
    .C1(_04336_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01834_));
 sky130_fd_sc_hd__mux2_1 _07765_ (.A0(\top.hTree.tree_reg[44] ),
    .A1(\top.findLeastValue.sum[44] ),
    .S(net286),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04338_));
 sky130_fd_sc_hd__mux2_1 _07766_ (.A0(\top.findLeastValue.sum[44] ),
    .A1(_04338_),
    .S(net392),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04339_));
 sky130_fd_sc_hd__or2_1 _07767_ (.A(net478),
    .B(_04338_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04340_));
 sky130_fd_sc_hd__o211a_1 _07768_ (.A1(net421),
    .A2(_04339_),
    .B1(_04340_),
    .C1(net262),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04341_));
 sky130_fd_sc_hd__a221o_1 _07769_ (.A1(net437),
    .A2(net1450),
    .B1(net252),
    .B2(\top.findLeastValue.sum[44] ),
    .C1(_04341_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01833_));
 sky130_fd_sc_hd__mux2_1 _07770_ (.A0(\top.hTree.tree_reg[43] ),
    .A1(\top.findLeastValue.sum[43] ),
    .S(net285),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04342_));
 sky130_fd_sc_hd__mux2_1 _07771_ (.A0(\top.hTree.tree_reg[43] ),
    .A1(\top.findLeastValue.sum[43] ),
    .S(_04251_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04343_));
 sky130_fd_sc_hd__or2_1 _07772_ (.A(net479),
    .B(_04342_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04344_));
 sky130_fd_sc_hd__o211a_1 _07773_ (.A1(net422),
    .A2(_04343_),
    .B1(_04344_),
    .C1(net262),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04345_));
 sky130_fd_sc_hd__a221o_1 _07774_ (.A1(net437),
    .A2(net1497),
    .B1(net252),
    .B2(\top.findLeastValue.sum[43] ),
    .C1(_04345_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01832_));
 sky130_fd_sc_hd__mux2_1 _07775_ (.A0(\top.hTree.tree_reg[42] ),
    .A1(\top.findLeastValue.sum[42] ),
    .S(net285),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04346_));
 sky130_fd_sc_hd__mux2_1 _07776_ (.A0(\top.hTree.tree_reg[42] ),
    .A1(\top.findLeastValue.sum[42] ),
    .S(net266),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04347_));
 sky130_fd_sc_hd__or2_1 _07777_ (.A(net479),
    .B(_04346_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04348_));
 sky130_fd_sc_hd__o211a_1 _07778_ (.A1(net420),
    .A2(_04347_),
    .B1(_04348_),
    .C1(net262),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04349_));
 sky130_fd_sc_hd__a221o_1 _07779_ (.A1(net437),
    .A2(net1569),
    .B1(net251),
    .B2(\top.findLeastValue.sum[42] ),
    .C1(_04349_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01831_));
 sky130_fd_sc_hd__mux2_1 _07780_ (.A0(\top.hTree.tree_reg[41] ),
    .A1(\top.findLeastValue.sum[41] ),
    .S(net285),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04350_));
 sky130_fd_sc_hd__mux2_1 _07781_ (.A0(\top.hTree.tree_reg[41] ),
    .A1(\top.findLeastValue.sum[41] ),
    .S(_04251_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04351_));
 sky130_fd_sc_hd__or2_1 _07782_ (.A(net479),
    .B(_04350_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04352_));
 sky130_fd_sc_hd__o211a_1 _07783_ (.A1(net420),
    .A2(_04351_),
    .B1(_04352_),
    .C1(net262),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04353_));
 sky130_fd_sc_hd__a221o_1 _07784_ (.A1(net437),
    .A2(net1645),
    .B1(net251),
    .B2(\top.findLeastValue.sum[41] ),
    .C1(_04353_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01830_));
 sky130_fd_sc_hd__mux2_1 _07785_ (.A0(\top.hTree.tree_reg[40] ),
    .A1(\top.findLeastValue.sum[40] ),
    .S(net285),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04354_));
 sky130_fd_sc_hd__mux2_1 _07786_ (.A0(\top.hTree.tree_reg[40] ),
    .A1(\top.findLeastValue.sum[40] ),
    .S(net267),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04355_));
 sky130_fd_sc_hd__or2_1 _07787_ (.A(net479),
    .B(_04354_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04356_));
 sky130_fd_sc_hd__o211a_1 _07788_ (.A1(net420),
    .A2(_04355_),
    .B1(_04356_),
    .C1(net262),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04357_));
 sky130_fd_sc_hd__a221o_1 _07789_ (.A1(net437),
    .A2(net1535),
    .B1(net251),
    .B2(\top.findLeastValue.sum[40] ),
    .C1(_04357_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01829_));
 sky130_fd_sc_hd__mux2_1 _07790_ (.A0(\top.hTree.tree_reg[39] ),
    .A1(\top.findLeastValue.sum[39] ),
    .S(net283),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04358_));
 sky130_fd_sc_hd__mux2_1 _07791_ (.A0(\top.hTree.tree_reg[39] ),
    .A1(\top.findLeastValue.sum[39] ),
    .S(net266),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04359_));
 sky130_fd_sc_hd__or2_1 _07792_ (.A(net476),
    .B(_04358_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04360_));
 sky130_fd_sc_hd__o211a_1 _07793_ (.A1(net418),
    .A2(_04359_),
    .B1(_04360_),
    .C1(net260),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04361_));
 sky130_fd_sc_hd__a221o_1 _07794_ (.A1(net435),
    .A2(net1610),
    .B1(net249),
    .B2(\top.findLeastValue.sum[39] ),
    .C1(_04361_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01828_));
 sky130_fd_sc_hd__mux2_1 _07795_ (.A0(\top.hTree.tree_reg[38] ),
    .A1(\top.findLeastValue.sum[38] ),
    .S(net283),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04362_));
 sky130_fd_sc_hd__mux2_1 _07796_ (.A0(\top.hTree.tree_reg[38] ),
    .A1(\top.findLeastValue.sum[38] ),
    .S(net266),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04363_));
 sky130_fd_sc_hd__or2_1 _07797_ (.A(net476),
    .B(_04362_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04364_));
 sky130_fd_sc_hd__o211a_1 _07798_ (.A1(net421),
    .A2(_04363_),
    .B1(_04364_),
    .C1(net260),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04365_));
 sky130_fd_sc_hd__a221o_1 _07799_ (.A1(net435),
    .A2(net1607),
    .B1(net252),
    .B2(\top.findLeastValue.sum[38] ),
    .C1(_04365_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01827_));
 sky130_fd_sc_hd__mux2_1 _07800_ (.A0(\top.hTree.tree_reg[37] ),
    .A1(\top.findLeastValue.sum[37] ),
    .S(net283),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04366_));
 sky130_fd_sc_hd__mux2_1 _07801_ (.A0(\top.hTree.tree_reg[37] ),
    .A1(\top.findLeastValue.sum[37] ),
    .S(net266),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04367_));
 sky130_fd_sc_hd__or2_1 _07802_ (.A(net476),
    .B(_04366_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04368_));
 sky130_fd_sc_hd__o211a_1 _07803_ (.A1(net418),
    .A2(_04367_),
    .B1(_04368_),
    .C1(net260),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04369_));
 sky130_fd_sc_hd__a221o_1 _07804_ (.A1(net435),
    .A2(net1594),
    .B1(net249),
    .B2(\top.findLeastValue.sum[37] ),
    .C1(_04369_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01826_));
 sky130_fd_sc_hd__mux2_1 _07805_ (.A0(\top.hTree.tree_reg[36] ),
    .A1(\top.findLeastValue.sum[36] ),
    .S(net283),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04370_));
 sky130_fd_sc_hd__mux2_1 _07806_ (.A0(\top.findLeastValue.sum[36] ),
    .A1(_04370_),
    .S(net391),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04371_));
 sky130_fd_sc_hd__or2_1 _07807_ (.A(net476),
    .B(_04370_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04372_));
 sky130_fd_sc_hd__o211a_1 _07808_ (.A1(net418),
    .A2(_04371_),
    .B1(_04372_),
    .C1(net260),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04373_));
 sky130_fd_sc_hd__a221o_1 _07809_ (.A1(net435),
    .A2(net1457),
    .B1(net249),
    .B2(\top.findLeastValue.sum[36] ),
    .C1(_04373_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01825_));
 sky130_fd_sc_hd__mux2_1 _07810_ (.A0(\top.hTree.tree_reg[35] ),
    .A1(\top.findLeastValue.sum[35] ),
    .S(net283),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04374_));
 sky130_fd_sc_hd__mux2_1 _07811_ (.A0(\top.findLeastValue.sum[35] ),
    .A1(_04374_),
    .S(net391),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04375_));
 sky130_fd_sc_hd__or2_1 _07812_ (.A(net476),
    .B(_04374_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04376_));
 sky130_fd_sc_hd__o211a_1 _07813_ (.A1(net418),
    .A2(_04375_),
    .B1(_04376_),
    .C1(net260),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04377_));
 sky130_fd_sc_hd__a221o_1 _07814_ (.A1(net435),
    .A2(net1492),
    .B1(net249),
    .B2(\top.findLeastValue.sum[35] ),
    .C1(_04377_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01824_));
 sky130_fd_sc_hd__mux2_1 _07815_ (.A0(\top.hTree.tree_reg[34] ),
    .A1(\top.findLeastValue.sum[34] ),
    .S(net283),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04378_));
 sky130_fd_sc_hd__mux2_1 _07816_ (.A0(\top.findLeastValue.sum[34] ),
    .A1(_04378_),
    .S(net391),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04379_));
 sky130_fd_sc_hd__or2_1 _07817_ (.A(net476),
    .B(_04378_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04380_));
 sky130_fd_sc_hd__o211a_1 _07818_ (.A1(net418),
    .A2(_04379_),
    .B1(_04380_),
    .C1(net260),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04381_));
 sky130_fd_sc_hd__a221o_1 _07819_ (.A1(net435),
    .A2(net1313),
    .B1(net249),
    .B2(\top.findLeastValue.sum[34] ),
    .C1(_04381_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01823_));
 sky130_fd_sc_hd__mux2_1 _07820_ (.A0(\top.hTree.tree_reg[33] ),
    .A1(\top.findLeastValue.sum[33] ),
    .S(net283),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04382_));
 sky130_fd_sc_hd__mux2_1 _07821_ (.A0(\top.hTree.tree_reg[33] ),
    .A1(\top.findLeastValue.sum[33] ),
    .S(net266),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04383_));
 sky130_fd_sc_hd__or2_1 _07822_ (.A(net476),
    .B(_04382_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04384_));
 sky130_fd_sc_hd__o211a_1 _07823_ (.A1(net418),
    .A2(_04383_),
    .B1(_04384_),
    .C1(net260),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04385_));
 sky130_fd_sc_hd__a221o_1 _07824_ (.A1(net435),
    .A2(net1585),
    .B1(net249),
    .B2(\top.findLeastValue.sum[33] ),
    .C1(_04385_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01822_));
 sky130_fd_sc_hd__mux2_1 _07825_ (.A0(\top.hTree.tree_reg[32] ),
    .A1(\top.findLeastValue.sum[32] ),
    .S(net283),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04386_));
 sky130_fd_sc_hd__mux2_1 _07826_ (.A0(\top.findLeastValue.sum[32] ),
    .A1(_04386_),
    .S(net391),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04387_));
 sky130_fd_sc_hd__or2_1 _07827_ (.A(net476),
    .B(_04386_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04388_));
 sky130_fd_sc_hd__o211a_1 _07828_ (.A1(net418),
    .A2(_04387_),
    .B1(_04388_),
    .C1(net260),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04389_));
 sky130_fd_sc_hd__a221o_1 _07829_ (.A1(net435),
    .A2(net1356),
    .B1(net249),
    .B2(\top.findLeastValue.sum[32] ),
    .C1(_04389_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01821_));
 sky130_fd_sc_hd__mux2_1 _07830_ (.A0(\top.hTree.tree_reg[31] ),
    .A1(\top.findLeastValue.sum[31] ),
    .S(net282),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04390_));
 sky130_fd_sc_hd__mux2_1 _07831_ (.A0(\top.hTree.tree_reg[31] ),
    .A1(\top.findLeastValue.sum[31] ),
    .S(net265),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04391_));
 sky130_fd_sc_hd__or2_1 _07832_ (.A(net470),
    .B(_04390_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04392_));
 sky130_fd_sc_hd__o211a_1 _07833_ (.A1(net417),
    .A2(_04391_),
    .B1(_04392_),
    .C1(net255),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04393_));
 sky130_fd_sc_hd__a221o_1 _07834_ (.A1(net431),
    .A2(net1537),
    .B1(net248),
    .B2(\top.findLeastValue.sum[31] ),
    .C1(_04393_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01820_));
 sky130_fd_sc_hd__mux2_1 _07835_ (.A0(\top.hTree.tree_reg[30] ),
    .A1(\top.findLeastValue.sum[30] ),
    .S(net282),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04394_));
 sky130_fd_sc_hd__mux2_1 _07836_ (.A0(\top.findLeastValue.sum[30] ),
    .A1(_04394_),
    .S(net390),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04395_));
 sky130_fd_sc_hd__or2_1 _07837_ (.A(net470),
    .B(_04394_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04396_));
 sky130_fd_sc_hd__o211a_1 _07838_ (.A1(net417),
    .A2(_04395_),
    .B1(_04396_),
    .C1(net255),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04397_));
 sky130_fd_sc_hd__a221o_1 _07839_ (.A1(net431),
    .A2(net1490),
    .B1(net248),
    .B2(\top.findLeastValue.sum[30] ),
    .C1(_04397_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01819_));
 sky130_fd_sc_hd__mux2_1 _07840_ (.A0(\top.hTree.tree_reg[29] ),
    .A1(\top.findLeastValue.sum[29] ),
    .S(net282),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04398_));
 sky130_fd_sc_hd__mux2_1 _07841_ (.A0(\top.findLeastValue.sum[29] ),
    .A1(_04398_),
    .S(net390),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04399_));
 sky130_fd_sc_hd__or2_1 _07842_ (.A(net470),
    .B(_04398_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04400_));
 sky130_fd_sc_hd__o211a_1 _07843_ (.A1(net417),
    .A2(_04399_),
    .B1(_04400_),
    .C1(net255),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04401_));
 sky130_fd_sc_hd__a221o_1 _07844_ (.A1(net434),
    .A2(net1493),
    .B1(net248),
    .B2(\top.findLeastValue.sum[29] ),
    .C1(_04401_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01818_));
 sky130_fd_sc_hd__mux2_1 _07845_ (.A0(\top.hTree.tree_reg[28] ),
    .A1(\top.findLeastValue.sum[28] ),
    .S(net282),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04402_));
 sky130_fd_sc_hd__mux2_1 _07846_ (.A0(\top.findLeastValue.sum[28] ),
    .A1(_04402_),
    .S(net390),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04403_));
 sky130_fd_sc_hd__or2_1 _07847_ (.A(net471),
    .B(_04402_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04404_));
 sky130_fd_sc_hd__o211a_1 _07848_ (.A1(net417),
    .A2(_04403_),
    .B1(_04404_),
    .C1(net256),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04405_));
 sky130_fd_sc_hd__a221o_1 _07849_ (.A1(net434),
    .A2(net1495),
    .B1(net248),
    .B2(net1801),
    .C1(_04405_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01817_));
 sky130_fd_sc_hd__mux2_1 _07850_ (.A0(\top.hTree.tree_reg[27] ),
    .A1(\top.findLeastValue.sum[27] ),
    .S(net282),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04406_));
 sky130_fd_sc_hd__mux2_1 _07851_ (.A0(\top.hTree.tree_reg[27] ),
    .A1(\top.findLeastValue.sum[27] ),
    .S(net265),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04407_));
 sky130_fd_sc_hd__or2_1 _07852_ (.A(net471),
    .B(_04406_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04408_));
 sky130_fd_sc_hd__o211a_1 _07853_ (.A1(net417),
    .A2(_04407_),
    .B1(_04408_),
    .C1(net259),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04409_));
 sky130_fd_sc_hd__a221o_1 _07854_ (.A1(net434),
    .A2(net1558),
    .B1(net248),
    .B2(\top.findLeastValue.sum[27] ),
    .C1(_04409_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01816_));
 sky130_fd_sc_hd__mux2_1 _07855_ (.A0(\top.hTree.tree_reg[26] ),
    .A1(\top.findLeastValue.sum[26] ),
    .S(net281),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04410_));
 sky130_fd_sc_hd__mux2_1 _07856_ (.A0(\top.hTree.tree_reg[26] ),
    .A1(\top.findLeastValue.sum[26] ),
    .S(net265),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04411_));
 sky130_fd_sc_hd__or2_1 _07857_ (.A(net475),
    .B(_04410_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04412_));
 sky130_fd_sc_hd__o211a_1 _07858_ (.A1(net422),
    .A2(_04411_),
    .B1(_04412_),
    .C1(net258),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04413_));
 sky130_fd_sc_hd__a221o_1 _07859_ (.A1(net432),
    .A2(net1546),
    .B1(net253),
    .B2(\top.findLeastValue.sum[26] ),
    .C1(_04413_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01815_));
 sky130_fd_sc_hd__mux2_1 _07860_ (.A0(\top.hTree.tree_reg[25] ),
    .A1(\top.findLeastValue.sum[25] ),
    .S(net281),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04414_));
 sky130_fd_sc_hd__mux2_1 _07861_ (.A0(\top.hTree.tree_reg[25] ),
    .A1(\top.findLeastValue.sum[25] ),
    .S(net264),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04415_));
 sky130_fd_sc_hd__or2_1 _07862_ (.A(net475),
    .B(_04414_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04416_));
 sky130_fd_sc_hd__o211a_1 _07863_ (.A1(net417),
    .A2(_04415_),
    .B1(_04416_),
    .C1(net258),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04417_));
 sky130_fd_sc_hd__a221o_1 _07864_ (.A1(net432),
    .A2(net1565),
    .B1(net253),
    .B2(\top.findLeastValue.sum[25] ),
    .C1(_04417_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01814_));
 sky130_fd_sc_hd__mux2_1 _07865_ (.A0(\top.hTree.tree_reg[24] ),
    .A1(\top.findLeastValue.sum[24] ),
    .S(net282),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04418_));
 sky130_fd_sc_hd__mux2_1 _07866_ (.A0(\top.findLeastValue.sum[24] ),
    .A1(_04418_),
    .S(net390),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04419_));
 sky130_fd_sc_hd__or2_1 _07867_ (.A(net471),
    .B(_04418_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04420_));
 sky130_fd_sc_hd__o211a_1 _07868_ (.A1(net422),
    .A2(_04419_),
    .B1(_04420_),
    .C1(net259),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04421_));
 sky130_fd_sc_hd__a221o_1 _07869_ (.A1(net431),
    .A2(net1431),
    .B1(net253),
    .B2(\top.findLeastValue.sum[24] ),
    .C1(_04421_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01813_));
 sky130_fd_sc_hd__mux2_1 _07870_ (.A0(\top.hTree.tree_reg[23] ),
    .A1(\top.findLeastValue.sum[23] ),
    .S(net281),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04422_));
 sky130_fd_sc_hd__mux2_1 _07871_ (.A0(\top.hTree.tree_reg[23] ),
    .A1(\top.findLeastValue.sum[23] ),
    .S(net264),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04423_));
 sky130_fd_sc_hd__or2_1 _07872_ (.A(net475),
    .B(_04422_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04424_));
 sky130_fd_sc_hd__o211a_1 _07873_ (.A1(net417),
    .A2(_04423_),
    .B1(_04424_),
    .C1(net258),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04425_));
 sky130_fd_sc_hd__a221o_1 _07874_ (.A1(net438),
    .A2(net1551),
    .B1(net248),
    .B2(net1806),
    .C1(_04425_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01812_));
 sky130_fd_sc_hd__mux2_1 _07875_ (.A0(\top.hTree.tree_reg[22] ),
    .A1(\top.findLeastValue.sum[22] ),
    .S(net281),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04426_));
 sky130_fd_sc_hd__mux2_1 _07876_ (.A0(\top.hTree.tree_reg[22] ),
    .A1(\top.findLeastValue.sum[22] ),
    .S(net265),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04427_));
 sky130_fd_sc_hd__or2_1 _07877_ (.A(net475),
    .B(_04426_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04428_));
 sky130_fd_sc_hd__o211a_1 _07878_ (.A1(net417),
    .A2(_04427_),
    .B1(_04428_),
    .C1(net263),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04429_));
 sky130_fd_sc_hd__a221o_1 _07879_ (.A1(net438),
    .A2(net1557),
    .B1(net248),
    .B2(net1807),
    .C1(_04429_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01811_));
 sky130_fd_sc_hd__mux2_1 _07880_ (.A0(\top.hTree.tree_reg[21] ),
    .A1(\top.findLeastValue.sum[21] ),
    .S(net281),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04430_));
 sky130_fd_sc_hd__mux2_1 _07881_ (.A0(\top.hTree.tree_reg[21] ),
    .A1(\top.findLeastValue.sum[21] ),
    .S(net264),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04431_));
 sky130_fd_sc_hd__or2_1 _07882_ (.A(net478),
    .B(_04430_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04432_));
 sky130_fd_sc_hd__o211a_1 _07883_ (.A1(net421),
    .A2(_04431_),
    .B1(_04432_),
    .C1(net263),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04433_));
 sky130_fd_sc_hd__a221o_1 _07884_ (.A1(net438),
    .A2(net1552),
    .B1(net248),
    .B2(\top.findLeastValue.sum[21] ),
    .C1(_04433_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01810_));
 sky130_fd_sc_hd__mux2_1 _07885_ (.A0(\top.hTree.tree_reg[20] ),
    .A1(\top.findLeastValue.sum[20] ),
    .S(net283),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04434_));
 sky130_fd_sc_hd__mux2_1 _07886_ (.A0(\top.findLeastValue.sum[20] ),
    .A1(_04434_),
    .S(net391),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04435_));
 sky130_fd_sc_hd__or2_1 _07887_ (.A(net476),
    .B(_04434_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04436_));
 sky130_fd_sc_hd__o211a_1 _07888_ (.A1(net421),
    .A2(_04435_),
    .B1(_04436_),
    .C1(net260),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04437_));
 sky130_fd_sc_hd__a221o_1 _07889_ (.A1(net435),
    .A2(net1395),
    .B1(net248),
    .B2(\top.findLeastValue.sum[20] ),
    .C1(_04437_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01809_));
 sky130_fd_sc_hd__mux2_1 _07890_ (.A0(\top.hTree.tree_reg[19] ),
    .A1(\top.findLeastValue.sum[19] ),
    .S(net286),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04438_));
 sky130_fd_sc_hd__mux2_1 _07891_ (.A0(\top.findLeastValue.sum[19] ),
    .A1(_04438_),
    .S(net392),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04439_));
 sky130_fd_sc_hd__or2_1 _07892_ (.A(net478),
    .B(_04438_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04440_));
 sky130_fd_sc_hd__o211a_1 _07893_ (.A1(net421),
    .A2(_04439_),
    .B1(_04440_),
    .C1(net263),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04441_));
 sky130_fd_sc_hd__a221o_1 _07894_ (.A1(net438),
    .A2(net1350),
    .B1(net252),
    .B2(\top.findLeastValue.sum[19] ),
    .C1(_04441_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01808_));
 sky130_fd_sc_hd__mux2_1 _07895_ (.A0(\top.hTree.tree_reg[18] ),
    .A1(\top.findLeastValue.sum[18] ),
    .S(net286),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04442_));
 sky130_fd_sc_hd__mux2_1 _07896_ (.A0(\top.hTree.tree_reg[18] ),
    .A1(\top.findLeastValue.sum[18] ),
    .S(net267),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04443_));
 sky130_fd_sc_hd__or2_1 _07897_ (.A(net478),
    .B(_04442_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04444_));
 sky130_fd_sc_hd__o211a_1 _07898_ (.A1(net421),
    .A2(_04443_),
    .B1(_04444_),
    .C1(net263),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04445_));
 sky130_fd_sc_hd__a221o_1 _07899_ (.A1(net438),
    .A2(net1570),
    .B1(net252),
    .B2(\top.findLeastValue.sum[18] ),
    .C1(_04445_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01807_));
 sky130_fd_sc_hd__mux2_1 _07900_ (.A0(\top.hTree.tree_reg[17] ),
    .A1(\top.findLeastValue.sum[17] ),
    .S(net286),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04446_));
 sky130_fd_sc_hd__mux2_1 _07901_ (.A0(\top.findLeastValue.sum[17] ),
    .A1(_04446_),
    .S(net392),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04447_));
 sky130_fd_sc_hd__or2_1 _07902_ (.A(net478),
    .B(_04446_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04448_));
 sky130_fd_sc_hd__o211a_1 _07903_ (.A1(net421),
    .A2(_04447_),
    .B1(_04448_),
    .C1(net263),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04449_));
 sky130_fd_sc_hd__a221o_1 _07904_ (.A1(net438),
    .A2(net1443),
    .B1(net252),
    .B2(\top.findLeastValue.sum[17] ),
    .C1(_04449_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01806_));
 sky130_fd_sc_hd__mux2_1 _07905_ (.A0(\top.hTree.tree_reg[16] ),
    .A1(\top.findLeastValue.sum[16] ),
    .S(net286),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04450_));
 sky130_fd_sc_hd__mux2_1 _07906_ (.A0(\top.hTree.tree_reg[16] ),
    .A1(\top.findLeastValue.sum[16] ),
    .S(net267),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04451_));
 sky130_fd_sc_hd__or2_1 _07907_ (.A(net478),
    .B(_04450_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04452_));
 sky130_fd_sc_hd__o211a_1 _07908_ (.A1(net421),
    .A2(_04451_),
    .B1(_04452_),
    .C1(net263),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04453_));
 sky130_fd_sc_hd__a221o_1 _07909_ (.A1(net438),
    .A2(net1567),
    .B1(net252),
    .B2(\top.findLeastValue.sum[16] ),
    .C1(_04453_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01805_));
 sky130_fd_sc_hd__mux2_1 _07910_ (.A0(\top.hTree.tree_reg[15] ),
    .A1(\top.findLeastValue.sum[15] ),
    .S(net286),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04454_));
 sky130_fd_sc_hd__mux2_1 _07911_ (.A0(\top.findLeastValue.sum[15] ),
    .A1(_04454_),
    .S(net391),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04455_));
 sky130_fd_sc_hd__or2_1 _07912_ (.A(net479),
    .B(_04454_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04456_));
 sky130_fd_sc_hd__o211a_1 _07913_ (.A1(net420),
    .A2(_04455_),
    .B1(_04456_),
    .C1(net262),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04457_));
 sky130_fd_sc_hd__a221o_1 _07914_ (.A1(net437),
    .A2(net1436),
    .B1(net251),
    .B2(\top.findLeastValue.sum[15] ),
    .C1(_04457_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01804_));
 sky130_fd_sc_hd__mux2_1 _07915_ (.A0(\top.hTree.tree_reg[14] ),
    .A1(\top.findLeastValue.sum[14] ),
    .S(net285),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04458_));
 sky130_fd_sc_hd__mux2_1 _07916_ (.A0(\top.hTree.tree_reg[14] ),
    .A1(\top.findLeastValue.sum[14] ),
    .S(net267),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04459_));
 sky130_fd_sc_hd__or2_1 _07917_ (.A(net479),
    .B(_04458_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04460_));
 sky130_fd_sc_hd__o211a_1 _07918_ (.A1(net420),
    .A2(_04459_),
    .B1(_04460_),
    .C1(net262),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04461_));
 sky130_fd_sc_hd__a221o_1 _07919_ (.A1(net437),
    .A2(net1584),
    .B1(net251),
    .B2(\top.findLeastValue.sum[14] ),
    .C1(_04461_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01803_));
 sky130_fd_sc_hd__mux2_1 _07920_ (.A0(\top.hTree.tree_reg[13] ),
    .A1(\top.findLeastValue.sum[13] ),
    .S(net285),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04462_));
 sky130_fd_sc_hd__mux2_1 _07921_ (.A0(\top.hTree.tree_reg[13] ),
    .A1(\top.findLeastValue.sum[13] ),
    .S(net267),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04463_));
 sky130_fd_sc_hd__or2_1 _07922_ (.A(net478),
    .B(_04462_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04464_));
 sky130_fd_sc_hd__o211a_1 _07923_ (.A1(net420),
    .A2(_04463_),
    .B1(_04464_),
    .C1(net262),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04465_));
 sky130_fd_sc_hd__a221o_1 _07924_ (.A1(net438),
    .A2(\top.hTree.tree_reg[13] ),
    .B1(net251),
    .B2(net1559),
    .C1(_04465_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01802_));
 sky130_fd_sc_hd__mux2_1 _07925_ (.A0(\top.hTree.tree_reg[12] ),
    .A1(\top.findLeastValue.sum[12] ),
    .S(net285),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04466_));
 sky130_fd_sc_hd__mux2_1 _07926_ (.A0(\top.findLeastValue.sum[12] ),
    .A1(_04466_),
    .S(net392),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04467_));
 sky130_fd_sc_hd__or2_1 _07927_ (.A(net478),
    .B(_04466_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04468_));
 sky130_fd_sc_hd__o211a_1 _07928_ (.A1(net420),
    .A2(_04467_),
    .B1(_04468_),
    .C1(net263),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04469_));
 sky130_fd_sc_hd__a221o_1 _07929_ (.A1(net437),
    .A2(net1433),
    .B1(net252),
    .B2(\top.findLeastValue.sum[12] ),
    .C1(_04469_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01801_));
 sky130_fd_sc_hd__mux2_1 _07930_ (.A0(\top.hTree.tree_reg[11] ),
    .A1(\top.findLeastValue.sum[11] ),
    .S(net285),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04470_));
 sky130_fd_sc_hd__mux2_1 _07931_ (.A0(\top.hTree.tree_reg[11] ),
    .A1(\top.findLeastValue.sum[11] ),
    .S(net267),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04471_));
 sky130_fd_sc_hd__or2_1 _07932_ (.A(net479),
    .B(_04470_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04472_));
 sky130_fd_sc_hd__o211a_1 _07933_ (.A1(net420),
    .A2(_04471_),
    .B1(_04472_),
    .C1(net262),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04473_));
 sky130_fd_sc_hd__a221o_1 _07934_ (.A1(net437),
    .A2(net1600),
    .B1(net251),
    .B2(\top.findLeastValue.sum[11] ),
    .C1(_04473_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01800_));
 sky130_fd_sc_hd__mux2_1 _07935_ (.A0(\top.hTree.tree_reg[10] ),
    .A1(\top.findLeastValue.sum[10] ),
    .S(net283),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04474_));
 sky130_fd_sc_hd__mux2_1 _07936_ (.A0(\top.hTree.tree_reg[10] ),
    .A1(\top.findLeastValue.sum[10] ),
    .S(net266),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04475_));
 sky130_fd_sc_hd__or2_1 _07937_ (.A(net477),
    .B(_04474_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04476_));
 sky130_fd_sc_hd__o211a_1 _07938_ (.A1(net418),
    .A2(_04475_),
    .B1(_04476_),
    .C1(net261),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04477_));
 sky130_fd_sc_hd__a221o_1 _07939_ (.A1(net436),
    .A2(net1589),
    .B1(net251),
    .B2(\top.findLeastValue.sum[10] ),
    .C1(_04477_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01799_));
 sky130_fd_sc_hd__mux2_1 _07940_ (.A0(\top.hTree.tree_reg[9] ),
    .A1(\top.findLeastValue.sum[9] ),
    .S(net285),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04478_));
 sky130_fd_sc_hd__mux2_1 _07941_ (.A0(\top.hTree.tree_reg[9] ),
    .A1(\top.findLeastValue.sum[9] ),
    .S(net266),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04479_));
 sky130_fd_sc_hd__or2_1 _07942_ (.A(net476),
    .B(_04478_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04480_));
 sky130_fd_sc_hd__o211a_1 _07943_ (.A1(net420),
    .A2(_04479_),
    .B1(_04480_),
    .C1(net260),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04481_));
 sky130_fd_sc_hd__a221o_1 _07944_ (.A1(net435),
    .A2(net1599),
    .B1(net251),
    .B2(\top.findLeastValue.sum[9] ),
    .C1(_04481_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01798_));
 sky130_fd_sc_hd__mux2_1 _07945_ (.A0(\top.hTree.tree_reg[8] ),
    .A1(\top.findLeastValue.sum[8] ),
    .S(net285),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04482_));
 sky130_fd_sc_hd__mux2_1 _07946_ (.A0(\top.hTree.tree_reg[8] ),
    .A1(\top.findLeastValue.sum[8] ),
    .S(net267),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04483_));
 sky130_fd_sc_hd__or2_1 _07947_ (.A(net478),
    .B(_04482_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04484_));
 sky130_fd_sc_hd__o211a_1 _07948_ (.A1(net420),
    .A2(_04483_),
    .B1(_04484_),
    .C1(net262),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04485_));
 sky130_fd_sc_hd__a221o_1 _07949_ (.A1(net437),
    .A2(net1564),
    .B1(net251),
    .B2(\top.findLeastValue.sum[8] ),
    .C1(_04485_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01797_));
 sky130_fd_sc_hd__mux2_1 _07950_ (.A0(\top.hTree.tree_reg[7] ),
    .A1(\top.findLeastValue.sum[7] ),
    .S(net284),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04486_));
 sky130_fd_sc_hd__mux2_1 _07951_ (.A0(\top.hTree.tree_reg[7] ),
    .A1(\top.findLeastValue.sum[7] ),
    .S(net266),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04487_));
 sky130_fd_sc_hd__or2_1 _07952_ (.A(net477),
    .B(_04486_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04488_));
 sky130_fd_sc_hd__o211a_1 _07953_ (.A1(net418),
    .A2(_04487_),
    .B1(_04488_),
    .C1(net261),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04489_));
 sky130_fd_sc_hd__a221o_1 _07954_ (.A1(net436),
    .A2(net1603),
    .B1(net249),
    .B2(net1800),
    .C1(_04489_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01796_));
 sky130_fd_sc_hd__mux2_1 _07955_ (.A0(\top.hTree.tree_reg[6] ),
    .A1(\top.findLeastValue.sum[6] ),
    .S(net284),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04490_));
 sky130_fd_sc_hd__mux2_1 _07956_ (.A0(\top.hTree.tree_reg[6] ),
    .A1(\top.findLeastValue.sum[6] ),
    .S(net266),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04491_));
 sky130_fd_sc_hd__or2_1 _07957_ (.A(net477),
    .B(_04490_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04492_));
 sky130_fd_sc_hd__o211a_1 _07958_ (.A1(net418),
    .A2(_04491_),
    .B1(_04492_),
    .C1(net261),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04493_));
 sky130_fd_sc_hd__a221o_1 _07959_ (.A1(net436),
    .A2(net1573),
    .B1(net250),
    .B2(\top.findLeastValue.sum[6] ),
    .C1(_04493_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01795_));
 sky130_fd_sc_hd__mux2_1 _07960_ (.A0(\top.hTree.tree_reg[5] ),
    .A1(\top.findLeastValue.sum[5] ),
    .S(net284),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04494_));
 sky130_fd_sc_hd__mux2_1 _07961_ (.A0(\top.hTree.tree_reg[5] ),
    .A1(\top.findLeastValue.sum[5] ),
    .S(net266),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04495_));
 sky130_fd_sc_hd__or2_1 _07962_ (.A(net477),
    .B(_04494_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04496_));
 sky130_fd_sc_hd__o211a_1 _07963_ (.A1(net419),
    .A2(_04495_),
    .B1(_04496_),
    .C1(net261),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04497_));
 sky130_fd_sc_hd__a221o_1 _07964_ (.A1(net436),
    .A2(net1579),
    .B1(net249),
    .B2(\top.findLeastValue.sum[5] ),
    .C1(_04497_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01794_));
 sky130_fd_sc_hd__mux2_1 _07965_ (.A0(\top.hTree.tree_reg[4] ),
    .A1(\top.findLeastValue.sum[4] ),
    .S(net284),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04498_));
 sky130_fd_sc_hd__mux2_1 _07966_ (.A0(\top.findLeastValue.sum[4] ),
    .A1(_04498_),
    .S(net391),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04499_));
 sky130_fd_sc_hd__or2_1 _07967_ (.A(net477),
    .B(_04498_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04500_));
 sky130_fd_sc_hd__o211a_1 _07968_ (.A1(net419),
    .A2(_04499_),
    .B1(_04500_),
    .C1(net261),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04501_));
 sky130_fd_sc_hd__a221o_1 _07969_ (.A1(net436),
    .A2(net1318),
    .B1(net249),
    .B2(\top.findLeastValue.sum[4] ),
    .C1(_04501_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01793_));
 sky130_fd_sc_hd__mux2_1 _07970_ (.A0(\top.hTree.tree_reg[3] ),
    .A1(\top.findLeastValue.sum[3] ),
    .S(net284),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04502_));
 sky130_fd_sc_hd__mux2_1 _07971_ (.A0(\top.findLeastValue.sum[3] ),
    .A1(_04502_),
    .S(net391),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04503_));
 sky130_fd_sc_hd__or2_1 _07972_ (.A(net477),
    .B(_04502_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04504_));
 sky130_fd_sc_hd__o211a_1 _07973_ (.A1(net419),
    .A2(_04503_),
    .B1(_04504_),
    .C1(net261),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04505_));
 sky130_fd_sc_hd__a221o_1 _07974_ (.A1(net436),
    .A2(net1229),
    .B1(net250),
    .B2(\top.findLeastValue.sum[3] ),
    .C1(_04505_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01792_));
 sky130_fd_sc_hd__mux2_1 _07975_ (.A0(\top.hTree.tree_reg[2] ),
    .A1(\top.findLeastValue.sum[2] ),
    .S(net284),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04506_));
 sky130_fd_sc_hd__mux2_1 _07976_ (.A0(\top.findLeastValue.sum[2] ),
    .A1(_04506_),
    .S(net391),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04507_));
 sky130_fd_sc_hd__or2_1 _07977_ (.A(net477),
    .B(_04506_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04508_));
 sky130_fd_sc_hd__o211a_1 _07978_ (.A1(net419),
    .A2(_04507_),
    .B1(_04508_),
    .C1(net261),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04509_));
 sky130_fd_sc_hd__a221o_1 _07979_ (.A1(net436),
    .A2(net1474),
    .B1(net250),
    .B2(\top.findLeastValue.sum[2] ),
    .C1(_04509_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01791_));
 sky130_fd_sc_hd__mux2_1 _07980_ (.A0(\top.hTree.tree_reg[1] ),
    .A1(\top.findLeastValue.sum[1] ),
    .S(net284),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04510_));
 sky130_fd_sc_hd__mux2_1 _07981_ (.A0(\top.hTree.tree_reg[1] ),
    .A1(\top.findLeastValue.sum[1] ),
    .S(net267),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04511_));
 sky130_fd_sc_hd__or2_1 _07982_ (.A(net477),
    .B(_04510_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04512_));
 sky130_fd_sc_hd__o211a_1 _07983_ (.A1(net419),
    .A2(_04511_),
    .B1(_04512_),
    .C1(net261),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04513_));
 sky130_fd_sc_hd__a221o_1 _07984_ (.A1(net436),
    .A2(net1538),
    .B1(net250),
    .B2(\top.findLeastValue.sum[1] ),
    .C1(_04513_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01790_));
 sky130_fd_sc_hd__mux2_1 _07985_ (.A0(\top.hTree.tree_reg[0] ),
    .A1(\top.findLeastValue.sum[0] ),
    .S(net284),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04514_));
 sky130_fd_sc_hd__mux2_1 _07986_ (.A0(\top.findLeastValue.sum[0] ),
    .A1(_04514_),
    .S(net391),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04515_));
 sky130_fd_sc_hd__or2_1 _07987_ (.A(net477),
    .B(_04514_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04516_));
 sky130_fd_sc_hd__o211a_1 _07988_ (.A1(net419),
    .A2(_04515_),
    .B1(_04516_),
    .C1(net261),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04517_));
 sky130_fd_sc_hd__a221o_1 _07989_ (.A1(net436),
    .A2(net1458),
    .B1(net250),
    .B2(\top.findLeastValue.sum[0] ),
    .C1(_04517_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01789_));
 sky130_fd_sc_hd__o21ai_1 _07990_ (.A1(\top.hTree.state[4] ),
    .A2(\top.hTree.state[3] ),
    .B1(net255),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04518_));
 sky130_fd_sc_hd__or2_1 _07991_ (.A(\top.hTree.state[5] ),
    .B(\top.hTree.state[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04519_));
 sky130_fd_sc_hd__o31a_1 _07992_ (.A1(\top.hTree.state[4] ),
    .A2(\top.hTree.state[3] ),
    .A3(_04519_),
    .B1(net254),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04520_));
 sky130_fd_sc_hd__a21o_1 _07993_ (.A1(net431),
    .A2(\top.WorR ),
    .B1(_04520_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01788_));
 sky130_fd_sc_hd__o21a_1 _07994_ (.A1(net448),
    .A2(net977),
    .B1(_04257_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01787_));
 sky130_fd_sc_hd__a21oi_1 _07995_ (.A1(\top.hTree.state[1] ),
    .A2(net254),
    .B1(net953),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04521_));
 sky130_fd_sc_hd__a21oi_1 _07996_ (.A1(net1004),
    .A2(net254),
    .B1(_04521_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_01786_));
 sky130_fd_sc_hd__o21a_2 _07997_ (.A1(_02846_),
    .A2(_04257_),
    .B1(_04518_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04522_));
 sky130_fd_sc_hd__nor2_2 _07998_ (.A(\top.hTree.state[6] ),
    .B(\top.hTree.state[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04523_));
 sky130_fd_sc_hd__mux2_1 _07999_ (.A0(\top.findLeastValue.least2[6] ),
    .A1(\top.findLeastValue.least1[6] ),
    .S(_04523_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04524_));
 sky130_fd_sc_hd__mux2_1 _08000_ (.A0(_04524_),
    .A1(net1728),
    .S(_04522_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01785_));
 sky130_fd_sc_hd__mux2_1 _08001_ (.A0(\top.findLeastValue.least2[5] ),
    .A1(\top.findLeastValue.least1[5] ),
    .S(_04523_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04525_));
 sky130_fd_sc_hd__mux2_1 _08002_ (.A0(_04525_),
    .A1(net1670),
    .S(_04522_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01784_));
 sky130_fd_sc_hd__mux2_1 _08003_ (.A0(\top.findLeastValue.least2[4] ),
    .A1(\top.findLeastValue.least1[4] ),
    .S(_04523_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04526_));
 sky130_fd_sc_hd__mux2_1 _08004_ (.A0(_04526_),
    .A1(net1695),
    .S(_04522_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01783_));
 sky130_fd_sc_hd__mux2_1 _08005_ (.A0(\top.findLeastValue.least2[3] ),
    .A1(\top.findLeastValue.least1[3] ),
    .S(_04523_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04527_));
 sky130_fd_sc_hd__mux2_1 _08006_ (.A0(_04527_),
    .A1(net1655),
    .S(_04522_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01782_));
 sky130_fd_sc_hd__mux2_1 _08007_ (.A0(\top.findLeastValue.least2[2] ),
    .A1(\top.findLeastValue.least1[2] ),
    .S(_04523_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04528_));
 sky130_fd_sc_hd__mux2_1 _08008_ (.A0(_04528_),
    .A1(net1618),
    .S(_04522_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01781_));
 sky130_fd_sc_hd__mux2_1 _08009_ (.A0(\top.findLeastValue.least2[1] ),
    .A1(\top.findLeastValue.least1[1] ),
    .S(_04523_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04529_));
 sky130_fd_sc_hd__mux2_1 _08010_ (.A0(_04529_),
    .A1(net1657),
    .S(_04522_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01780_));
 sky130_fd_sc_hd__mux2_1 _08011_ (.A0(\top.findLeastValue.least2[0] ),
    .A1(\top.findLeastValue.least1[0] ),
    .S(_04523_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04530_));
 sky130_fd_sc_hd__mux2_1 _08012_ (.A0(_04530_),
    .A1(net1672),
    .S(_04522_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01779_));
 sky130_fd_sc_hd__a22o_1 _08013_ (.A1(net1699),
    .A2(_04518_),
    .B1(_04519_),
    .B2(net254),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01778_));
 sky130_fd_sc_hd__nand2_1 _08014_ (.A(\top.findLeastValue.alternator_timer[1] ),
    .B(\top.findLeastValue.alternator_timer[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04531_));
 sky130_fd_sc_hd__a41o_1 _08015_ (.A1(\top.findLeastValue.alternator_timer[2] ),
    .A2(\top.findLeastValue.alternator_timer[1] ),
    .A3(\top.findLeastValue.alternator_timer[0] ),
    .A4(_03666_),
    .B1(\top.findLeastValue.alternator_timer[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04532_));
 sky130_fd_sc_hd__nor2_1 _08016_ (.A(net406),
    .B(_02790_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04533_));
 sky130_fd_sc_hd__o211a_1 _08017_ (.A1(_02562_),
    .A2(_04533_),
    .B1(_04532_),
    .C1(net287),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01777_));
 sky130_fd_sc_hd__a31o_1 _08018_ (.A1(\top.findLeastValue.alternator_timer[1] ),
    .A2(\top.findLeastValue.alternator_timer[0] ),
    .A3(_03666_),
    .B1(\top.findLeastValue.alternator_timer[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04534_));
 sky130_fd_sc_hd__a21oi_1 _08019_ (.A1(\top.findLeastValue.alternator_timer[2] ),
    .A2(net406),
    .B1(_02790_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04535_));
 sky130_fd_sc_hd__nand2_1 _08020_ (.A(_02783_),
    .B(_04535_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04536_));
 sky130_fd_sc_hd__a32o_1 _08021_ (.A1(\top.findLeastValue.alternator_timer[2] ),
    .A2(\top.findLeastValue.alternator_timer[1] ),
    .A3(\top.findLeastValue.alternator_timer[0] ),
    .B1(_02785_),
    .B2(_04536_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04537_));
 sky130_fd_sc_hd__nand2_1 _08022_ (.A(net456),
    .B(_04537_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04538_));
 sky130_fd_sc_hd__and3_1 _08023_ (.A(net287),
    .B(_04534_),
    .C(_04538_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01776_));
 sky130_fd_sc_hd__and3_1 _08024_ (.A(_02784_),
    .B(_03395_),
    .C(_04531_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04539_));
 sky130_fd_sc_hd__a22o_1 _08025_ (.A1(\top.findLeastValue.alternator_timer[1] ),
    .A2(_03665_),
    .B1(_04535_),
    .B2(_04539_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01775_));
 sky130_fd_sc_hd__nor2_1 _08026_ (.A(\top.findLeastValue.alternator_timer[0] ),
    .B(_02791_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04540_));
 sky130_fd_sc_hd__a22o_1 _08027_ (.A1(\top.findLeastValue.alternator_timer[0] ),
    .A2(_03665_),
    .B1(_04540_),
    .B2(_03395_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01774_));
 sky130_fd_sc_hd__nand2_1 _08028_ (.A(net514),
    .B(net463),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04541_));
 sky130_fd_sc_hd__nor2_1 _08029_ (.A(\top.CB_write_complete ),
    .B(_04541_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04542_));
 sky130_fd_sc_hd__nand2_1 _08030_ (.A(\top.CB_read_complete ),
    .B(\top.cb_syn.setup ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04543_));
 sky130_fd_sc_hd__and3_1 _08031_ (.A(\top.CB_read_complete ),
    .B(\top.cb_syn.setup ),
    .C(_04542_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04544_));
 sky130_fd_sc_hd__nor2_1 _08032_ (.A(_02525_),
    .B(_04544_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_01773_));
 sky130_fd_sc_hd__or3_1 _08033_ (.A(net514),
    .B(\top.cb_syn.curr_state[0] ),
    .C(_04181_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04545_));
 sky130_fd_sc_hd__nand2_1 _08034_ (.A(\top.cb_syn.setup ),
    .B(net463),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04546_));
 sky130_fd_sc_hd__and3_1 _08035_ (.A(\top.cb_syn.setup ),
    .B(net463),
    .C(\top.cb_syn.curr_state[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04547_));
 sky130_fd_sc_hd__nand2b_1 _08036_ (.A_N(\top.cb_syn.end_cond ),
    .B(\top.CB_write_complete ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04548_));
 sky130_fd_sc_hd__a21o_1 _08037_ (.A1(net514),
    .A2(_04548_),
    .B1(net423),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04549_));
 sky130_fd_sc_hd__and4bb_1 _08038_ (.A_N(_04549_),
    .B_N(_04547_),
    .C(_04545_),
    .D(_02891_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04550_));
 sky130_fd_sc_hd__nor2_1 _08039_ (.A(net550),
    .B(_02580_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04551_));
 sky130_fd_sc_hd__or4b_1 _08040_ (.A(net488),
    .B(net550),
    .C(net412),
    .D_N(net524),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04552_));
 sky130_fd_sc_hd__nand2_1 _08041_ (.A(net550),
    .B(_02894_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04553_));
 sky130_fd_sc_hd__and3_1 _08042_ (.A(net524),
    .B(_02889_),
    .C(_04553_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04554_));
 sky130_fd_sc_hd__or4_1 _08043_ (.A(net515),
    .B(net514),
    .C(_02886_),
    .D(_04554_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04555_));
 sky130_fd_sc_hd__mux2_1 _08044_ (.A0(net488),
    .A1(_04555_),
    .S(_04550_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01772_));
 sky130_fd_sc_hd__a21oi_1 _08045_ (.A1(net550),
    .A2(_04189_),
    .B1(_04188_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04556_));
 sky130_fd_sc_hd__nor2_1 _08046_ (.A(_04190_),
    .B(_04556_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04557_));
 sky130_fd_sc_hd__a211o_1 _08047_ (.A1(net523),
    .A2(_02995_),
    .B1(_04204_),
    .C1(_04557_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04558_));
 sky130_fd_sc_hd__inv_2 _08048_ (.A(_04558_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04559_));
 sky130_fd_sc_hd__and2_1 _08049_ (.A(net523),
    .B(_02969_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04560_));
 sky130_fd_sc_hd__nor2_1 _08050_ (.A(_04207_),
    .B(_04560_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04561_));
 sky130_fd_sc_hd__and2_1 _08051_ (.A(\top.cb_syn.char_path_n[1] ),
    .B(_04201_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04562_));
 sky130_fd_sc_hd__nand2_1 _08052_ (.A(\top.cb_syn.char_path_n[2] ),
    .B(_04562_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04563_));
 sky130_fd_sc_hd__o41a_1 _08053_ (.A1(net515),
    .A2(net522),
    .A3(net523),
    .A4(net514),
    .B1(_04561_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04564_));
 sky130_fd_sc_hd__a21bo_1 _08054_ (.A1(net515),
    .A2(_04563_),
    .B1_N(_04564_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04565_));
 sky130_fd_sc_hd__a211o_2 _08055_ (.A1(net514),
    .A2(_04548_),
    .B1(_04558_),
    .C1(_04565_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04566_));
 sky130_fd_sc_hd__nand2_1 _08056_ (.A(\top.cb_syn.zeroes[1] ),
    .B(\top.cb_syn.zeroes[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04567_));
 sky130_fd_sc_hd__or2_1 _08057_ (.A(_02531_),
    .B(_04567_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04568_));
 sky130_fd_sc_hd__nor2_1 _08058_ (.A(_02530_),
    .B(_04568_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04569_));
 sky130_fd_sc_hd__inv_2 _08059_ (.A(_04569_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04570_));
 sky130_fd_sc_hd__nand2_1 _08060_ (.A(\top.cb_syn.zeroes[4] ),
    .B(_04569_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04571_));
 sky130_fd_sc_hd__nor2_1 _08061_ (.A(_02528_),
    .B(_04571_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04572_));
 sky130_fd_sc_hd__inv_2 _08062_ (.A(_04572_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04573_));
 sky130_fd_sc_hd__nand2_1 _08063_ (.A(\top.cb_syn.zeroes[6] ),
    .B(_04572_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04574_));
 sky130_fd_sc_hd__a21o_1 _08064_ (.A1(_04179_),
    .A2(_04574_),
    .B1(_04566_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04575_));
 sky130_fd_sc_hd__and2b_2 _08065_ (.A_N(_04566_),
    .B(_04179_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04576_));
 sky130_fd_sc_hd__nor2_1 _08066_ (.A(\top.cb_syn.zeroes[7] ),
    .B(_04574_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04577_));
 sky130_fd_sc_hd__a22o_1 _08067_ (.A1(\top.cb_syn.zeroes[7] ),
    .A2(_04575_),
    .B1(_04576_),
    .B2(_04577_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01771_));
 sky130_fd_sc_hd__nor2_1 _08068_ (.A(_04566_),
    .B(_04573_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04578_));
 sky130_fd_sc_hd__o21a_1 _08069_ (.A1(net1726),
    .A2(_04578_),
    .B1(_04575_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01770_));
 sky130_fd_sc_hd__nand2_1 _08070_ (.A(_02528_),
    .B(_04571_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04579_));
 sky130_fd_sc_hd__a32o_1 _08071_ (.A1(_04573_),
    .A2(_04576_),
    .A3(_04579_),
    .B1(_04566_),
    .B2(\top.cb_syn.zeroes[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01769_));
 sky130_fd_sc_hd__or2_1 _08072_ (.A(\top.cb_syn.zeroes[4] ),
    .B(_04569_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04580_));
 sky130_fd_sc_hd__a32o_1 _08073_ (.A1(_04571_),
    .A2(_04576_),
    .A3(_04580_),
    .B1(_04566_),
    .B2(net1787),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01768_));
 sky130_fd_sc_hd__nand2_1 _08074_ (.A(_02530_),
    .B(_04568_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04581_));
 sky130_fd_sc_hd__a32o_1 _08075_ (.A1(_04570_),
    .A2(_04576_),
    .A3(_04581_),
    .B1(_04566_),
    .B2(net1722),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01767_));
 sky130_fd_sc_hd__nand2_1 _08076_ (.A(_02531_),
    .B(_04567_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04582_));
 sky130_fd_sc_hd__a32o_1 _08077_ (.A1(_04568_),
    .A2(_04576_),
    .A3(_04582_),
    .B1(_04566_),
    .B2(net1703),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01766_));
 sky130_fd_sc_hd__a32o_1 _08078_ (.A1(_03386_),
    .A2(_04567_),
    .A3(_04576_),
    .B1(_04566_),
    .B2(net1717),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01765_));
 sky130_fd_sc_hd__mux2_1 _08079_ (.A0(_04566_),
    .A1(_04576_),
    .S(_02533_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01764_));
 sky130_fd_sc_hd__o21a_1 _08080_ (.A1(net550),
    .A2(_02890_),
    .B1(net524),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04583_));
 sky130_fd_sc_hd__nor2_1 _08081_ (.A(_04549_),
    .B(_04552_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04584_));
 sky130_fd_sc_hd__o32a_1 _08082_ (.A1(_04541_),
    .A2(_04548_),
    .A3(_04583_),
    .B1(_04584_),
    .B2(net1085),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01763_));
 sky130_fd_sc_hd__nor2_1 _08083_ (.A(_04203_),
    .B(_04551_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04585_));
 sky130_fd_sc_hd__a2bb2o_1 _08084_ (.A1_N(\top.cb_syn.check_right ),
    .A2_N(_04552_),
    .B1(_02896_),
    .B2(net412),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04586_));
 sky130_fd_sc_hd__a211o_1 _08085_ (.A1(net488),
    .A2(_04178_),
    .B1(_04585_),
    .C1(_04586_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04587_));
 sky130_fd_sc_hd__or3_1 _08086_ (.A(net519),
    .B(net524),
    .C(net514),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04588_));
 sky130_fd_sc_hd__or4b_4 _08087_ (.A(_04196_),
    .B(_04549_),
    .C(_04587_),
    .D_N(_04588_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04589_));
 sky130_fd_sc_hd__nor3_4 _08088_ (.A(net519),
    .B(net514),
    .C(_04589_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04590_));
 sky130_fd_sc_hd__nand2_1 _08089_ (.A(\top.cb_syn.num_lefts[1] ),
    .B(\top.cb_syn.num_lefts[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04591_));
 sky130_fd_sc_hd__and3_1 _08090_ (.A(\top.cb_syn.num_lefts[2] ),
    .B(\top.cb_syn.num_lefts[1] ),
    .C(\top.cb_syn.num_lefts[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04592_));
 sky130_fd_sc_hd__inv_2 _08091_ (.A(_04592_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04593_));
 sky130_fd_sc_hd__nand2_1 _08092_ (.A(\top.cb_syn.num_lefts[3] ),
    .B(_04592_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04594_));
 sky130_fd_sc_hd__and4_1 _08093_ (.A(\top.cb_syn.num_lefts[5] ),
    .B(\top.cb_syn.num_lefts[4] ),
    .C(\top.cb_syn.num_lefts[3] ),
    .D(_04592_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04595_));
 sky130_fd_sc_hd__inv_2 _08094_ (.A(_04595_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04596_));
 sky130_fd_sc_hd__nand2_1 _08095_ (.A(\top.cb_syn.num_lefts[6] ),
    .B(_04595_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04597_));
 sky130_fd_sc_hd__xnor2_1 _08096_ (.A(\top.cb_syn.num_lefts[7] ),
    .B(_04597_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04598_));
 sky130_fd_sc_hd__a22o_1 _08097_ (.A1(\top.cb_syn.num_lefts[7] ),
    .A2(_04589_),
    .B1(_04590_),
    .B2(_04598_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01762_));
 sky130_fd_sc_hd__or2_1 _08098_ (.A(\top.cb_syn.num_lefts[6] ),
    .B(_04595_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04599_));
 sky130_fd_sc_hd__a32o_1 _08099_ (.A1(_04590_),
    .A2(_04597_),
    .A3(_04599_),
    .B1(_04589_),
    .B2(net1682),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01761_));
 sky130_fd_sc_hd__a31o_1 _08100_ (.A1(\top.cb_syn.num_lefts[4] ),
    .A2(\top.cb_syn.num_lefts[3] ),
    .A3(_04592_),
    .B1(\top.cb_syn.num_lefts[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04600_));
 sky130_fd_sc_hd__a32o_1 _08101_ (.A1(_04590_),
    .A2(_04596_),
    .A3(_04600_),
    .B1(_04589_),
    .B2(net1661),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01760_));
 sky130_fd_sc_hd__xnor2_1 _08102_ (.A(\top.cb_syn.num_lefts[4] ),
    .B(_04594_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04601_));
 sky130_fd_sc_hd__a22o_1 _08103_ (.A1(\top.cb_syn.num_lefts[4] ),
    .A2(_04589_),
    .B1(_04590_),
    .B2(_04601_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01759_));
 sky130_fd_sc_hd__or2_1 _08104_ (.A(\top.cb_syn.num_lefts[3] ),
    .B(_04592_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04602_));
 sky130_fd_sc_hd__a32o_1 _08105_ (.A1(_04590_),
    .A2(_04594_),
    .A3(_04602_),
    .B1(_04589_),
    .B2(\top.cb_syn.num_lefts[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01758_));
 sky130_fd_sc_hd__a21o_1 _08106_ (.A1(\top.cb_syn.num_lefts[1] ),
    .A2(\top.cb_syn.num_lefts[0] ),
    .B1(\top.cb_syn.num_lefts[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04603_));
 sky130_fd_sc_hd__a32o_1 _08107_ (.A1(_04590_),
    .A2(_04593_),
    .A3(_04603_),
    .B1(_04589_),
    .B2(net1660),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01757_));
 sky130_fd_sc_hd__or2_1 _08108_ (.A(\top.cb_syn.num_lefts[1] ),
    .B(\top.cb_syn.num_lefts[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04604_));
 sky130_fd_sc_hd__a32o_1 _08109_ (.A1(_04590_),
    .A2(_04591_),
    .A3(_04604_),
    .B1(_04589_),
    .B2(\top.cb_syn.num_lefts[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01756_));
 sky130_fd_sc_hd__mux2_1 _08110_ (.A0(_04590_),
    .A1(_04589_),
    .S(\top.cb_syn.num_lefts[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01755_));
 sky130_fd_sc_hd__and2_1 _08111_ (.A(net523),
    .B(_02994_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04605_));
 sky130_fd_sc_hd__nor2_1 _08112_ (.A(\top.cb_syn.h_element[54] ),
    .B(net412),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04606_));
 sky130_fd_sc_hd__or3_1 _08113_ (.A(net489),
    .B(_04195_),
    .C(_04606_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04607_));
 sky130_fd_sc_hd__nand2_1 _08114_ (.A(net464),
    .B(_04607_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04608_));
 sky130_fd_sc_hd__a221o_1 _08115_ (.A1(net412),
    .A2(_02887_),
    .B1(_04178_),
    .B2(net489),
    .C1(_04585_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04609_));
 sky130_fd_sc_hd__a311o_1 _08116_ (.A1(_02539_),
    .A2(_02886_),
    .A3(_04606_),
    .B1(_04608_),
    .C1(_04609_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04610_));
 sky130_fd_sc_hd__nor2_1 _08117_ (.A(net515),
    .B(\top.cb_syn.curr_state[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04611_));
 sky130_fd_sc_hd__or2_2 _08118_ (.A(net515),
    .B(net523),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04612_));
 sky130_fd_sc_hd__nor2_1 _08119_ (.A(_04178_),
    .B(net370),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04613_));
 sky130_fd_sc_hd__or4_1 _08120_ (.A(_04202_),
    .B(_04586_),
    .C(_04610_),
    .D(_04613_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04614_));
 sky130_fd_sc_hd__nor3_2 _08121_ (.A(_04560_),
    .B(_04605_),
    .C(_04614_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04615_));
 sky130_fd_sc_hd__or3_2 _08122_ (.A(_04560_),
    .B(_04605_),
    .C(_04614_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04616_));
 sky130_fd_sc_hd__and4_1 _08123_ (.A(\top.cb_syn.cb_length[2] ),
    .B(\top.cb_syn.cb_length[1] ),
    .C(\top.cb_syn.cb_length[0] ),
    .D(_04611_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04617_));
 sky130_fd_sc_hd__nand2_1 _08124_ (.A(\top.cb_syn.cb_length[3] ),
    .B(_04617_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04618_));
 sky130_fd_sc_hd__nor2_1 _08125_ (.A(_04200_),
    .B(_04611_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04619_));
 sky130_fd_sc_hd__nand2_1 _08126_ (.A(_02535_),
    .B(_04619_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04620_));
 sky130_fd_sc_hd__and2_1 _08127_ (.A(_02534_),
    .B(_04620_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04621_));
 sky130_fd_sc_hd__a211o_1 _08128_ (.A1(\top.cb_syn.cb_length[4] ),
    .A2(_04618_),
    .B1(_04621_),
    .C1(net172),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04622_));
 sky130_fd_sc_hd__nand2_1 _08129_ (.A(\top.cb_syn.cb_length[5] ),
    .B(_04611_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04623_));
 sky130_fd_sc_hd__or2_1 _08130_ (.A(\top.cb_syn.cb_length[5] ),
    .B(_04611_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04624_));
 sky130_fd_sc_hd__a21oi_1 _08131_ (.A1(_04623_),
    .A2(_04624_),
    .B1(_04622_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04625_));
 sky130_fd_sc_hd__xor2_1 _08132_ (.A(net1470),
    .B(_04625_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01754_));
 sky130_fd_sc_hd__xnor2_1 _08133_ (.A(net1723),
    .B(_04622_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_01753_));
 sky130_fd_sc_hd__a21oi_1 _08134_ (.A1(_04618_),
    .A2(_04620_),
    .B1(net172),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04626_));
 sky130_fd_sc_hd__xnor2_1 _08135_ (.A(_02534_),
    .B(_04626_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_01752_));
 sky130_fd_sc_hd__o21a_1 _08136_ (.A1(_04617_),
    .A2(_04619_),
    .B1(net190),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04627_));
 sky130_fd_sc_hd__xnor2_1 _08137_ (.A(_02535_),
    .B(_04627_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_01751_));
 sky130_fd_sc_hd__or2_1 _08138_ (.A(\top.cb_syn.cb_length[2] ),
    .B(net190),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04628_));
 sky130_fd_sc_hd__o21ai_1 _08139_ (.A1(\top.cb_syn.cb_length[1] ),
    .A2(\top.cb_syn.cb_length[0] ),
    .B1(\top.cb_syn.cb_length[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04629_));
 sky130_fd_sc_hd__nand2b_1 _08140_ (.A_N(\top.cb_syn.cb_length[1] ),
    .B(\top.cb_syn.cb_length[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04630_));
 sky130_fd_sc_hd__nand2b_1 _08141_ (.A_N(\top.cb_syn.cb_length[0] ),
    .B(\top.cb_syn.cb_length[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04631_));
 sky130_fd_sc_hd__and3_1 _08142_ (.A(_04611_),
    .B(_04630_),
    .C(_04631_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04632_));
 sky130_fd_sc_hd__and3_1 _08143_ (.A(_04200_),
    .B(_04629_),
    .C(_04632_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04633_));
 sky130_fd_sc_hd__a21oi_1 _08144_ (.A1(_04200_),
    .A2(_04629_),
    .B1(_04632_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04634_));
 sky130_fd_sc_hd__o31a_1 _08145_ (.A1(net172),
    .A2(_04633_),
    .A3(_04634_),
    .B1(_04628_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01750_));
 sky130_fd_sc_hd__a21oi_1 _08146_ (.A1(_04630_),
    .A2(_04631_),
    .B1(_04611_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04635_));
 sky130_fd_sc_hd__nor2_1 _08147_ (.A(_04632_),
    .B(_04635_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04636_));
 sky130_fd_sc_hd__mux2_1 _08148_ (.A0(\top.cb_syn.cb_length[1] ),
    .A1(_04636_),
    .S(net190),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01749_));
 sky130_fd_sc_hd__xnor2_1 _08149_ (.A(\top.cb_syn.cb_length[0] ),
    .B(net172),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_01748_));
 sky130_fd_sc_hd__nand2_1 _08150_ (.A(_02538_),
    .B(net371),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04637_));
 sky130_fd_sc_hd__and3_1 _08151_ (.A(\top.cb_syn.char_path_n[127] ),
    .B(net190),
    .C(net326),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04638_));
 sky130_fd_sc_hd__a21o_1 _08152_ (.A1(net1555),
    .A2(net172),
    .B1(_04638_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01747_));
 sky130_fd_sc_hd__a221o_1 _08153_ (.A1(\top.cb_syn.curr_path[127] ),
    .A2(net369),
    .B1(net326),
    .B2(\top.cb_syn.char_path_n[126] ),
    .C1(net172),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04639_));
 sky130_fd_sc_hd__o21a_1 _08154_ (.A1(\top.cb_syn.char_path_n[127] ),
    .A2(net190),
    .B1(_04639_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01746_));
 sky130_fd_sc_hd__a221o_1 _08155_ (.A1(\top.cb_syn.char_path_n[127] ),
    .A2(net370),
    .B1(net328),
    .B2(\top.cb_syn.char_path_n[125] ),
    .C1(net174),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04640_));
 sky130_fd_sc_hd__o21a_1 _08156_ (.A1(net1771),
    .A2(net192),
    .B1(_04640_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01745_));
 sky130_fd_sc_hd__a221o_1 _08157_ (.A1(\top.cb_syn.char_path_n[126] ),
    .A2(net370),
    .B1(net328),
    .B2(\top.cb_syn.char_path_n[124] ),
    .C1(net174),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04641_));
 sky130_fd_sc_hd__o21a_1 _08158_ (.A1(\top.cb_syn.char_path_n[125] ),
    .A2(net192),
    .B1(_04641_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01744_));
 sky130_fd_sc_hd__a221o_1 _08159_ (.A1(\top.cb_syn.char_path_n[125] ),
    .A2(net369),
    .B1(net326),
    .B2(\top.cb_syn.char_path_n[123] ),
    .C1(net173),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04642_));
 sky130_fd_sc_hd__o21a_1 _08160_ (.A1(net1785),
    .A2(net191),
    .B1(_04642_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01743_));
 sky130_fd_sc_hd__a221o_1 _08161_ (.A1(\top.cb_syn.char_path_n[124] ),
    .A2(net369),
    .B1(net326),
    .B2(\top.cb_syn.char_path_n[122] ),
    .C1(net173),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04643_));
 sky130_fd_sc_hd__o21a_1 _08162_ (.A1(\top.cb_syn.char_path_n[123] ),
    .A2(net191),
    .B1(_04643_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01742_));
 sky130_fd_sc_hd__a221o_1 _08163_ (.A1(\top.cb_syn.char_path_n[123] ),
    .A2(net369),
    .B1(net326),
    .B2(\top.cb_syn.char_path_n[121] ),
    .C1(net173),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04644_));
 sky130_fd_sc_hd__o21a_1 _08164_ (.A1(\top.cb_syn.char_path_n[122] ),
    .A2(net191),
    .B1(_04644_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01741_));
 sky130_fd_sc_hd__a221o_1 _08165_ (.A1(\top.cb_syn.char_path_n[122] ),
    .A2(net373),
    .B1(net327),
    .B2(\top.cb_syn.char_path_n[120] ),
    .C1(net176),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04645_));
 sky130_fd_sc_hd__o21a_1 _08166_ (.A1(\top.cb_syn.char_path_n[121] ),
    .A2(net194),
    .B1(_04645_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01740_));
 sky130_fd_sc_hd__a221o_1 _08167_ (.A1(\top.cb_syn.char_path_n[121] ),
    .A2(net373),
    .B1(net331),
    .B2(\top.cb_syn.char_path_n[119] ),
    .C1(net176),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04646_));
 sky130_fd_sc_hd__o21a_1 _08168_ (.A1(\top.cb_syn.char_path_n[120] ),
    .A2(net194),
    .B1(_04646_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01739_));
 sky130_fd_sc_hd__a221o_1 _08169_ (.A1(\top.cb_syn.char_path_n[120] ),
    .A2(net374),
    .B1(net330),
    .B2(\top.cb_syn.char_path_n[118] ),
    .C1(net177),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04647_));
 sky130_fd_sc_hd__o21a_1 _08170_ (.A1(net1738),
    .A2(net195),
    .B1(_04647_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01738_));
 sky130_fd_sc_hd__a221o_1 _08171_ (.A1(\top.cb_syn.char_path_n[119] ),
    .A2(net371),
    .B1(net329),
    .B2(\top.cb_syn.char_path_n[117] ),
    .C1(net175),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04648_));
 sky130_fd_sc_hd__o21a_1 _08172_ (.A1(\top.cb_syn.char_path_n[118] ),
    .A2(net193),
    .B1(_04648_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01737_));
 sky130_fd_sc_hd__a221o_1 _08173_ (.A1(\top.cb_syn.char_path_n[118] ),
    .A2(net377),
    .B1(net330),
    .B2(\top.cb_syn.char_path_n[116] ),
    .C1(net180),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04649_));
 sky130_fd_sc_hd__o21a_1 _08174_ (.A1(net1710),
    .A2(net198),
    .B1(_04649_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01736_));
 sky130_fd_sc_hd__a221o_1 _08175_ (.A1(\top.cb_syn.char_path_n[117] ),
    .A2(net377),
    .B1(net334),
    .B2(\top.cb_syn.char_path_n[115] ),
    .C1(net180),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04650_));
 sky130_fd_sc_hd__o21a_1 _08176_ (.A1(\top.cb_syn.char_path_n[116] ),
    .A2(net198),
    .B1(_04650_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01735_));
 sky130_fd_sc_hd__a221o_1 _08177_ (.A1(\top.cb_syn.char_path_n[116] ),
    .A2(net377),
    .B1(net334),
    .B2(\top.cb_syn.char_path_n[114] ),
    .C1(net180),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04651_));
 sky130_fd_sc_hd__o21a_1 _08178_ (.A1(\top.cb_syn.char_path_n[115] ),
    .A2(net198),
    .B1(_04651_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01734_));
 sky130_fd_sc_hd__a221o_1 _08179_ (.A1(\top.cb_syn.char_path_n[115] ),
    .A2(net378),
    .B1(net334),
    .B2(\top.cb_syn.char_path_n[113] ),
    .C1(net181),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04652_));
 sky130_fd_sc_hd__o21a_1 _08180_ (.A1(net1737),
    .A2(net199),
    .B1(_04652_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01733_));
 sky130_fd_sc_hd__a221o_1 _08181_ (.A1(\top.cb_syn.char_path_n[114] ),
    .A2(net378),
    .B1(net335),
    .B2(\top.cb_syn.char_path_n[112] ),
    .C1(net181),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04653_));
 sky130_fd_sc_hd__o21a_1 _08182_ (.A1(net1755),
    .A2(net199),
    .B1(_04653_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01732_));
 sky130_fd_sc_hd__a221o_1 _08183_ (.A1(\top.cb_syn.char_path_n[113] ),
    .A2(net378),
    .B1(net334),
    .B2(\top.cb_syn.char_path_n[111] ),
    .C1(net181),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04654_));
 sky130_fd_sc_hd__o21a_1 _08184_ (.A1(net1759),
    .A2(net199),
    .B1(_04654_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01731_));
 sky130_fd_sc_hd__a221o_1 _08185_ (.A1(\top.cb_syn.char_path_n[112] ),
    .A2(net385),
    .B1(net340),
    .B2(\top.cb_syn.char_path_n[110] ),
    .C1(net188),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04655_));
 sky130_fd_sc_hd__o21a_1 _08186_ (.A1(net1744),
    .A2(net205),
    .B1(_04655_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01730_));
 sky130_fd_sc_hd__a221o_1 _08187_ (.A1(\top.cb_syn.char_path_n[111] ),
    .A2(net383),
    .B1(net339),
    .B2(\top.cb_syn.char_path_n[109] ),
    .C1(net186),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04656_));
 sky130_fd_sc_hd__o21a_1 _08188_ (.A1(\top.cb_syn.char_path_n[110] ),
    .A2(net203),
    .B1(_04656_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01729_));
 sky130_fd_sc_hd__a221o_1 _08189_ (.A1(\top.cb_syn.char_path_n[110] ),
    .A2(net383),
    .B1(net339),
    .B2(\top.cb_syn.char_path_n[108] ),
    .C1(net186),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04657_));
 sky130_fd_sc_hd__o21a_1 _08190_ (.A1(\top.cb_syn.char_path_n[109] ),
    .A2(net203),
    .B1(_04657_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01728_));
 sky130_fd_sc_hd__a221o_1 _08191_ (.A1(\top.cb_syn.char_path_n[109] ),
    .A2(net383),
    .B1(net339),
    .B2(\top.cb_syn.char_path_n[107] ),
    .C1(net186),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04658_));
 sky130_fd_sc_hd__o21a_1 _08192_ (.A1(net1772),
    .A2(net203),
    .B1(_04658_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01727_));
 sky130_fd_sc_hd__a221o_1 _08193_ (.A1(\top.cb_syn.char_path_n[108] ),
    .A2(net383),
    .B1(net339),
    .B2(\top.cb_syn.char_path_n[106] ),
    .C1(net186),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04659_));
 sky130_fd_sc_hd__o21a_1 _08194_ (.A1(\top.cb_syn.char_path_n[107] ),
    .A2(net203),
    .B1(_04659_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01726_));
 sky130_fd_sc_hd__a221o_1 _08195_ (.A1(\top.cb_syn.char_path_n[107] ),
    .A2(net383),
    .B1(net339),
    .B2(\top.cb_syn.char_path_n[105] ),
    .C1(net186),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04660_));
 sky130_fd_sc_hd__o21a_1 _08196_ (.A1(\top.cb_syn.char_path_n[106] ),
    .A2(net203),
    .B1(_04660_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01725_));
 sky130_fd_sc_hd__a221o_1 _08197_ (.A1(\top.cb_syn.char_path_n[106] ),
    .A2(net381),
    .B1(net337),
    .B2(\top.cb_syn.char_path_n[104] ),
    .C1(net183),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04661_));
 sky130_fd_sc_hd__o21a_1 _08198_ (.A1(net1765),
    .A2(net201),
    .B1(_04661_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01724_));
 sky130_fd_sc_hd__a221o_1 _08199_ (.A1(\top.cb_syn.char_path_n[105] ),
    .A2(net380),
    .B1(net337),
    .B2(\top.cb_syn.char_path_n[103] ),
    .C1(net183),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04662_));
 sky130_fd_sc_hd__o21a_1 _08200_ (.A1(\top.cb_syn.char_path_n[104] ),
    .A2(net201),
    .B1(_04662_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01723_));
 sky130_fd_sc_hd__a221o_1 _08201_ (.A1(\top.cb_syn.char_path_n[104] ),
    .A2(net380),
    .B1(net337),
    .B2(\top.cb_syn.char_path_n[102] ),
    .C1(net183),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04663_));
 sky130_fd_sc_hd__o21a_1 _08202_ (.A1(\top.cb_syn.char_path_n[103] ),
    .A2(net201),
    .B1(_04663_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01722_));
 sky130_fd_sc_hd__a221o_1 _08203_ (.A1(\top.cb_syn.char_path_n[103] ),
    .A2(net380),
    .B1(net337),
    .B2(\top.cb_syn.char_path_n[101] ),
    .C1(net183),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04664_));
 sky130_fd_sc_hd__o21a_1 _08204_ (.A1(\top.cb_syn.char_path_n[102] ),
    .A2(net201),
    .B1(_04664_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01721_));
 sky130_fd_sc_hd__a221o_1 _08205_ (.A1(\top.cb_syn.char_path_n[102] ),
    .A2(net380),
    .B1(net336),
    .B2(\top.cb_syn.char_path_n[100] ),
    .C1(net183),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04665_));
 sky130_fd_sc_hd__o21a_1 _08206_ (.A1(\top.cb_syn.char_path_n[101] ),
    .A2(net201),
    .B1(_04665_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01720_));
 sky130_fd_sc_hd__a221o_1 _08207_ (.A1(\top.cb_syn.char_path_n[101] ),
    .A2(net379),
    .B1(net336),
    .B2(\top.cb_syn.char_path_n[99] ),
    .C1(net182),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04666_));
 sky130_fd_sc_hd__o21a_1 _08208_ (.A1(net1770),
    .A2(net200),
    .B1(_04666_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01719_));
 sky130_fd_sc_hd__a221o_1 _08209_ (.A1(\top.cb_syn.char_path_n[100] ),
    .A2(net379),
    .B1(net336),
    .B2(\top.cb_syn.char_path_n[98] ),
    .C1(net182),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04667_));
 sky130_fd_sc_hd__o21a_1 _08210_ (.A1(\top.cb_syn.char_path_n[99] ),
    .A2(net200),
    .B1(_04667_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01718_));
 sky130_fd_sc_hd__a221o_1 _08211_ (.A1(\top.cb_syn.char_path_n[99] ),
    .A2(net380),
    .B1(net336),
    .B2(\top.cb_syn.char_path_n[97] ),
    .C1(net183),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04668_));
 sky130_fd_sc_hd__o21a_1 _08212_ (.A1(\top.cb_syn.char_path_n[98] ),
    .A2(net200),
    .B1(_04668_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01717_));
 sky130_fd_sc_hd__a221o_1 _08213_ (.A1(\top.cb_syn.char_path_n[98] ),
    .A2(net372),
    .B1(net329),
    .B2(\top.cb_syn.char_path_n[96] ),
    .C1(net177),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04669_));
 sky130_fd_sc_hd__o21a_1 _08214_ (.A1(\top.cb_syn.char_path_n[97] ),
    .A2(net195),
    .B1(_04669_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01716_));
 sky130_fd_sc_hd__a221o_1 _08215_ (.A1(\top.cb_syn.char_path_n[97] ),
    .A2(net370),
    .B1(net328),
    .B2(\top.cb_syn.char_path_n[95] ),
    .C1(net174),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04670_));
 sky130_fd_sc_hd__o21a_1 _08216_ (.A1(\top.cb_syn.char_path_n[96] ),
    .A2(net192),
    .B1(_04670_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01715_));
 sky130_fd_sc_hd__a221o_1 _08217_ (.A1(\top.cb_syn.char_path_n[96] ),
    .A2(net370),
    .B1(net326),
    .B2(\top.cb_syn.char_path_n[94] ),
    .C1(net172),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04671_));
 sky130_fd_sc_hd__o21a_1 _08218_ (.A1(\top.cb_syn.char_path_n[95] ),
    .A2(net190),
    .B1(_04671_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01714_));
 sky130_fd_sc_hd__a221o_1 _08219_ (.A1(\top.cb_syn.char_path_n[95] ),
    .A2(net369),
    .B1(net326),
    .B2(\top.cb_syn.char_path_n[93] ),
    .C1(net173),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04672_));
 sky130_fd_sc_hd__o21a_1 _08220_ (.A1(net1794),
    .A2(net191),
    .B1(_04672_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01713_));
 sky130_fd_sc_hd__a221o_1 _08221_ (.A1(\top.cb_syn.char_path_n[94] ),
    .A2(net370),
    .B1(net326),
    .B2(\top.cb_syn.char_path_n[92] ),
    .C1(net172),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04673_));
 sky130_fd_sc_hd__o21a_1 _08222_ (.A1(\top.cb_syn.char_path_n[93] ),
    .A2(net191),
    .B1(_04673_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01712_));
 sky130_fd_sc_hd__a221o_1 _08223_ (.A1(\top.cb_syn.char_path_n[93] ),
    .A2(net369),
    .B1(net326),
    .B2(\top.cb_syn.char_path_n[91] ),
    .C1(net172),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04674_));
 sky130_fd_sc_hd__o21a_1 _08224_ (.A1(net1788),
    .A2(net190),
    .B1(_04674_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01711_));
 sky130_fd_sc_hd__a221o_1 _08225_ (.A1(\top.cb_syn.char_path_n[92] ),
    .A2(net369),
    .B1(net327),
    .B2(\top.cb_syn.char_path_n[90] ),
    .C1(net173),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04675_));
 sky130_fd_sc_hd__o21a_1 _08226_ (.A1(net1721),
    .A2(net190),
    .B1(_04675_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01710_));
 sky130_fd_sc_hd__a221o_1 _08227_ (.A1(\top.cb_syn.char_path_n[91] ),
    .A2(net369),
    .B1(net326),
    .B2(\top.cb_syn.char_path_n[89] ),
    .C1(net173),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04676_));
 sky130_fd_sc_hd__o21a_1 _08228_ (.A1(\top.cb_syn.char_path_n[90] ),
    .A2(net190),
    .B1(_04676_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01709_));
 sky130_fd_sc_hd__a221o_1 _08229_ (.A1(\top.cb_syn.char_path_n[90] ),
    .A2(net373),
    .B1(net331),
    .B2(\top.cb_syn.char_path_n[88] ),
    .C1(net176),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04677_));
 sky130_fd_sc_hd__o21a_1 _08230_ (.A1(net1746),
    .A2(net194),
    .B1(_04677_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01708_));
 sky130_fd_sc_hd__a221o_1 _08231_ (.A1(\top.cb_syn.char_path_n[89] ),
    .A2(net373),
    .B1(net327),
    .B2(\top.cb_syn.char_path_n[87] ),
    .C1(net176),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04678_));
 sky130_fd_sc_hd__o21a_1 _08232_ (.A1(\top.cb_syn.char_path_n[88] ),
    .A2(net194),
    .B1(_04678_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01707_));
 sky130_fd_sc_hd__a221o_1 _08233_ (.A1(\top.cb_syn.char_path_n[88] ),
    .A2(net377),
    .B1(net330),
    .B2(\top.cb_syn.char_path_n[86] ),
    .C1(net180),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04679_));
 sky130_fd_sc_hd__o21a_1 _08234_ (.A1(\top.cb_syn.char_path_n[87] ),
    .A2(net198),
    .B1(_04679_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01706_));
 sky130_fd_sc_hd__a221o_1 _08235_ (.A1(\top.cb_syn.char_path_n[87] ),
    .A2(net377),
    .B1(net334),
    .B2(\top.cb_syn.char_path_n[85] ),
    .C1(net180),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04680_));
 sky130_fd_sc_hd__o21a_1 _08236_ (.A1(\top.cb_syn.char_path_n[86] ),
    .A2(net198),
    .B1(_04680_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01705_));
 sky130_fd_sc_hd__a221o_1 _08237_ (.A1(\top.cb_syn.char_path_n[86] ),
    .A2(net377),
    .B1(net334),
    .B2(\top.cb_syn.char_path_n[84] ),
    .C1(net180),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04681_));
 sky130_fd_sc_hd__o21a_1 _08238_ (.A1(\top.cb_syn.char_path_n[85] ),
    .A2(net198),
    .B1(_04681_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01704_));
 sky130_fd_sc_hd__a221o_1 _08239_ (.A1(\top.cb_syn.char_path_n[85] ),
    .A2(net378),
    .B1(net334),
    .B2(\top.cb_syn.char_path_n[83] ),
    .C1(net180),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04682_));
 sky130_fd_sc_hd__o21a_1 _08240_ (.A1(net1767),
    .A2(net198),
    .B1(_04682_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01703_));
 sky130_fd_sc_hd__a221o_1 _08241_ (.A1(\top.cb_syn.char_path_n[84] ),
    .A2(net377),
    .B1(net334),
    .B2(\top.cb_syn.char_path_n[82] ),
    .C1(net180),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04683_));
 sky130_fd_sc_hd__o21a_1 _08242_ (.A1(net1720),
    .A2(net198),
    .B1(_04683_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01702_));
 sky130_fd_sc_hd__a221o_1 _08243_ (.A1(\top.cb_syn.char_path_n[83] ),
    .A2(net378),
    .B1(net335),
    .B2(\top.cb_syn.char_path_n[81] ),
    .C1(net181),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04684_));
 sky130_fd_sc_hd__o21a_1 _08244_ (.A1(net1752),
    .A2(net199),
    .B1(_04684_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01701_));
 sky130_fd_sc_hd__a221o_1 _08245_ (.A1(\top.cb_syn.char_path_n[82] ),
    .A2(net385),
    .B1(net335),
    .B2(\top.cb_syn.char_path_n[80] ),
    .C1(net188),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04685_));
 sky130_fd_sc_hd__o21a_1 _08246_ (.A1(net1736),
    .A2(net199),
    .B1(_04685_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01700_));
 sky130_fd_sc_hd__a221o_1 _08247_ (.A1(\top.cb_syn.char_path_n[81] ),
    .A2(net385),
    .B1(net340),
    .B2(\top.cb_syn.char_path_n[79] ),
    .C1(net188),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04686_));
 sky130_fd_sc_hd__o21a_1 _08248_ (.A1(net1719),
    .A2(net205),
    .B1(_04686_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01699_));
 sky130_fd_sc_hd__a221o_1 _08249_ (.A1(\top.cb_syn.char_path_n[80] ),
    .A2(net385),
    .B1(net340),
    .B2(\top.cb_syn.char_path_n[78] ),
    .C1(net188),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04687_));
 sky130_fd_sc_hd__o21a_1 _08250_ (.A1(\top.cb_syn.char_path_n[79] ),
    .A2(net205),
    .B1(_04687_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01698_));
 sky130_fd_sc_hd__a221o_1 _08251_ (.A1(\top.cb_syn.char_path_n[79] ),
    .A2(net384),
    .B1(net339),
    .B2(\top.cb_syn.char_path_n[77] ),
    .C1(net186),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04688_));
 sky130_fd_sc_hd__o21a_1 _08252_ (.A1(\top.cb_syn.char_path_n[78] ),
    .A2(net203),
    .B1(_04688_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01697_));
 sky130_fd_sc_hd__a221o_1 _08253_ (.A1(\top.cb_syn.char_path_n[78] ),
    .A2(net384),
    .B1(net339),
    .B2(\top.cb_syn.char_path_n[76] ),
    .C1(net187),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04689_));
 sky130_fd_sc_hd__o21a_1 _08254_ (.A1(\top.cb_syn.char_path_n[77] ),
    .A2(net204),
    .B1(_04689_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01696_));
 sky130_fd_sc_hd__a221o_1 _08255_ (.A1(\top.cb_syn.char_path_n[77] ),
    .A2(net384),
    .B1(net339),
    .B2(\top.cb_syn.char_path_n[75] ),
    .C1(net186),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04690_));
 sky130_fd_sc_hd__o21a_1 _08256_ (.A1(net1741),
    .A2(net203),
    .B1(_04690_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01695_));
 sky130_fd_sc_hd__a221o_1 _08257_ (.A1(\top.cb_syn.char_path_n[76] ),
    .A2(net383),
    .B1(net339),
    .B2(\top.cb_syn.char_path_n[74] ),
    .C1(net186),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04691_));
 sky130_fd_sc_hd__o21a_1 _08258_ (.A1(net1792),
    .A2(net203),
    .B1(_04691_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01694_));
 sky130_fd_sc_hd__a221o_1 _08259_ (.A1(\top.cb_syn.char_path_n[75] ),
    .A2(net383),
    .B1(net341),
    .B2(\top.cb_syn.char_path_n[73] ),
    .C1(net186),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04692_));
 sky130_fd_sc_hd__o21a_1 _08260_ (.A1(\top.cb_syn.char_path_n[74] ),
    .A2(net203),
    .B1(_04692_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01693_));
 sky130_fd_sc_hd__a221o_1 _08261_ (.A1(\top.cb_syn.char_path_n[74] ),
    .A2(net380),
    .B1(net337),
    .B2(\top.cb_syn.char_path_n[72] ),
    .C1(net183),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04693_));
 sky130_fd_sc_hd__o21a_1 _08262_ (.A1(\top.cb_syn.char_path_n[73] ),
    .A2(net201),
    .B1(_04693_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01692_));
 sky130_fd_sc_hd__a221o_1 _08263_ (.A1(\top.cb_syn.char_path_n[73] ),
    .A2(net380),
    .B1(net337),
    .B2(\top.cb_syn.char_path_n[71] ),
    .C1(net184),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04694_));
 sky130_fd_sc_hd__o21a_1 _08264_ (.A1(\top.cb_syn.char_path_n[72] ),
    .A2(net201),
    .B1(_04694_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01691_));
 sky130_fd_sc_hd__a221o_1 _08265_ (.A1(\top.cb_syn.char_path_n[72] ),
    .A2(net379),
    .B1(net336),
    .B2(\top.cb_syn.char_path_n[70] ),
    .C1(net182),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04695_));
 sky130_fd_sc_hd__o21a_1 _08266_ (.A1(\top.cb_syn.char_path_n[71] ),
    .A2(net202),
    .B1(_04695_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01690_));
 sky130_fd_sc_hd__a221o_1 _08267_ (.A1(\top.cb_syn.char_path_n[71] ),
    .A2(net376),
    .B1(net333),
    .B2(\top.cb_syn.char_path_n[69] ),
    .C1(net178),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04696_));
 sky130_fd_sc_hd__o21a_1 _08268_ (.A1(net1763),
    .A2(net196),
    .B1(_04696_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01689_));
 sky130_fd_sc_hd__a221o_1 _08269_ (.A1(\top.cb_syn.char_path_n[70] ),
    .A2(net375),
    .B1(net333),
    .B2(\top.cb_syn.char_path_n[68] ),
    .C1(net178),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04697_));
 sky130_fd_sc_hd__o21a_1 _08270_ (.A1(net1773),
    .A2(net196),
    .B1(_04697_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01688_));
 sky130_fd_sc_hd__a221o_1 _08271_ (.A1(\top.cb_syn.char_path_n[69] ),
    .A2(net375),
    .B1(net333),
    .B2(\top.cb_syn.char_path_n[67] ),
    .C1(net178),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04698_));
 sky130_fd_sc_hd__o21a_1 _08272_ (.A1(\top.cb_syn.char_path_n[68] ),
    .A2(net196),
    .B1(_04698_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01687_));
 sky130_fd_sc_hd__a221o_1 _08273_ (.A1(\top.cb_syn.char_path_n[68] ),
    .A2(net375),
    .B1(net333),
    .B2(\top.cb_syn.char_path_n[66] ),
    .C1(net178),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04699_));
 sky130_fd_sc_hd__o21a_1 _08274_ (.A1(\top.cb_syn.char_path_n[67] ),
    .A2(net196),
    .B1(_04699_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01686_));
 sky130_fd_sc_hd__a221o_1 _08275_ (.A1(\top.cb_syn.char_path_n[67] ),
    .A2(net375),
    .B1(net333),
    .B2(\top.cb_syn.char_path_n[65] ),
    .C1(net178),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04700_));
 sky130_fd_sc_hd__o21a_1 _08276_ (.A1(\top.cb_syn.char_path_n[66] ),
    .A2(net196),
    .B1(_04700_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01685_));
 sky130_fd_sc_hd__a221o_1 _08277_ (.A1(\top.cb_syn.char_path_n[66] ),
    .A2(net372),
    .B1(net329),
    .B2(\top.cb_syn.char_path_n[64] ),
    .C1(net177),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04701_));
 sky130_fd_sc_hd__o21a_1 _08278_ (.A1(\top.cb_syn.char_path_n[65] ),
    .A2(net195),
    .B1(_04701_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01684_));
 sky130_fd_sc_hd__a221o_1 _08279_ (.A1(\top.cb_syn.char_path_n[65] ),
    .A2(net372),
    .B1(net329),
    .B2(\top.cb_syn.char_path_n[63] ),
    .C1(net175),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04702_));
 sky130_fd_sc_hd__o21a_1 _08280_ (.A1(\top.cb_syn.char_path_n[64] ),
    .A2(net193),
    .B1(_04702_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01683_));
 sky130_fd_sc_hd__a221o_1 _08281_ (.A1(\top.cb_syn.char_path_n[64] ),
    .A2(net371),
    .B1(net328),
    .B2(\top.cb_syn.char_path_n[62] ),
    .C1(net175),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04703_));
 sky130_fd_sc_hd__o21a_1 _08282_ (.A1(net1745),
    .A2(net193),
    .B1(_04703_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01682_));
 sky130_fd_sc_hd__a221o_1 _08283_ (.A1(\top.cb_syn.char_path_n[63] ),
    .A2(net370),
    .B1(net328),
    .B2(\top.cb_syn.char_path_n[61] ),
    .C1(net174),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04704_));
 sky130_fd_sc_hd__o21a_1 _08284_ (.A1(\top.cb_syn.char_path_n[62] ),
    .A2(net192),
    .B1(_04704_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01681_));
 sky130_fd_sc_hd__a221o_1 _08285_ (.A1(\top.cb_syn.char_path_n[62] ),
    .A2(net371),
    .B1(net328),
    .B2(\top.cb_syn.char_path_n[60] ),
    .C1(net175),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04705_));
 sky130_fd_sc_hd__o21a_1 _08286_ (.A1(\top.cb_syn.char_path_n[61] ),
    .A2(net193),
    .B1(_04705_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01680_));
 sky130_fd_sc_hd__a221o_1 _08287_ (.A1(\top.cb_syn.char_path_n[61] ),
    .A2(net371),
    .B1(net328),
    .B2(\top.cb_syn.char_path_n[59] ),
    .C1(net174),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04706_));
 sky130_fd_sc_hd__o21a_1 _08288_ (.A1(\top.cb_syn.char_path_n[60] ),
    .A2(net192),
    .B1(_04706_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01679_));
 sky130_fd_sc_hd__a221o_1 _08289_ (.A1(\top.cb_syn.char_path_n[60] ),
    .A2(net371),
    .B1(net328),
    .B2(\top.cb_syn.char_path_n[58] ),
    .C1(net175),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04707_));
 sky130_fd_sc_hd__o21a_1 _08290_ (.A1(\top.cb_syn.char_path_n[59] ),
    .A2(net193),
    .B1(_04707_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01678_));
 sky130_fd_sc_hd__a221o_1 _08291_ (.A1(\top.cb_syn.char_path_n[59] ),
    .A2(net371),
    .B1(net328),
    .B2(\top.cb_syn.char_path_n[57] ),
    .C1(net175),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04708_));
 sky130_fd_sc_hd__o21a_1 _08292_ (.A1(\top.cb_syn.char_path_n[58] ),
    .A2(net193),
    .B1(_04708_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01677_));
 sky130_fd_sc_hd__a221o_1 _08293_ (.A1(\top.cb_syn.char_path_n[58] ),
    .A2(net371),
    .B1(net329),
    .B2(\top.cb_syn.char_path_n[56] ),
    .C1(net177),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04709_));
 sky130_fd_sc_hd__o21a_1 _08294_ (.A1(\top.cb_syn.char_path_n[57] ),
    .A2(net193),
    .B1(_04709_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01676_));
 sky130_fd_sc_hd__a221o_1 _08295_ (.A1(\top.cb_syn.char_path_n[57] ),
    .A2(net371),
    .B1(net329),
    .B2(\top.cb_syn.char_path_n[55] ),
    .C1(net175),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04710_));
 sky130_fd_sc_hd__o21a_1 _08296_ (.A1(\top.cb_syn.char_path_n[56] ),
    .A2(net195),
    .B1(_04710_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01675_));
 sky130_fd_sc_hd__a221o_1 _08297_ (.A1(\top.cb_syn.char_path_n[56] ),
    .A2(net372),
    .B1(net329),
    .B2(\top.cb_syn.char_path_n[54] ),
    .C1(net175),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04711_));
 sky130_fd_sc_hd__o21a_1 _08298_ (.A1(\top.cb_syn.char_path_n[55] ),
    .A2(net193),
    .B1(_04711_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01674_));
 sky130_fd_sc_hd__a221o_1 _08299_ (.A1(\top.cb_syn.char_path_n[55] ),
    .A2(net372),
    .B1(net329),
    .B2(\top.cb_syn.char_path_n[53] ),
    .C1(net175),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04712_));
 sky130_fd_sc_hd__o21a_1 _08300_ (.A1(\top.cb_syn.char_path_n[54] ),
    .A2(net193),
    .B1(_04712_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01673_));
 sky130_fd_sc_hd__a221o_1 _08301_ (.A1(\top.cb_syn.char_path_n[54] ),
    .A2(net376),
    .B1(net329),
    .B2(\top.cb_syn.char_path_n[52] ),
    .C1(net179),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04713_));
 sky130_fd_sc_hd__o21a_1 _08302_ (.A1(net1692),
    .A2(net197),
    .B1(_04713_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01672_));
 sky130_fd_sc_hd__a221o_1 _08303_ (.A1(\top.cb_syn.char_path_n[53] ),
    .A2(net376),
    .B1(net332),
    .B2(\top.cb_syn.char_path_n[51] ),
    .C1(net179),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04714_));
 sky130_fd_sc_hd__o21a_1 _08304_ (.A1(net1697),
    .A2(net197),
    .B1(_04714_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01671_));
 sky130_fd_sc_hd__a221o_1 _08305_ (.A1(\top.cb_syn.char_path_n[52] ),
    .A2(net376),
    .B1(net332),
    .B2(\top.cb_syn.char_path_n[50] ),
    .C1(net179),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04715_));
 sky130_fd_sc_hd__o21a_1 _08306_ (.A1(net1756),
    .A2(net197),
    .B1(_04715_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01670_));
 sky130_fd_sc_hd__a221o_1 _08307_ (.A1(\top.cb_syn.char_path_n[51] ),
    .A2(net375),
    .B1(net332),
    .B2(\top.cb_syn.char_path_n[49] ),
    .C1(net178),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04716_));
 sky130_fd_sc_hd__o21a_1 _08308_ (.A1(net1747),
    .A2(net196),
    .B1(_04716_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01669_));
 sky130_fd_sc_hd__a221o_1 _08309_ (.A1(\top.cb_syn.char_path_n[50] ),
    .A2(net376),
    .B1(net333),
    .B2(\top.cb_syn.char_path_n[48] ),
    .C1(net179),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04717_));
 sky130_fd_sc_hd__o21a_1 _08310_ (.A1(\top.cb_syn.char_path_n[49] ),
    .A2(net196),
    .B1(_04717_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01668_));
 sky130_fd_sc_hd__a221o_1 _08311_ (.A1(\top.cb_syn.char_path_n[49] ),
    .A2(net375),
    .B1(net333),
    .B2(\top.cb_syn.char_path_n[47] ),
    .C1(net178),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04718_));
 sky130_fd_sc_hd__o21a_1 _08312_ (.A1(\top.cb_syn.char_path_n[48] ),
    .A2(net196),
    .B1(_04718_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01667_));
 sky130_fd_sc_hd__a221o_1 _08313_ (.A1(\top.cb_syn.char_path_n[48] ),
    .A2(net382),
    .B1(net332),
    .B2(\top.cb_syn.char_path_n[46] ),
    .C1(net185),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04719_));
 sky130_fd_sc_hd__o21a_1 _08314_ (.A1(\top.cb_syn.char_path_n[47] ),
    .A2(net202),
    .B1(_04719_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01666_));
 sky130_fd_sc_hd__a221o_1 _08315_ (.A1(\top.cb_syn.char_path_n[47] ),
    .A2(net382),
    .B1(net338),
    .B2(\top.cb_syn.char_path_n[45] ),
    .C1(net185),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04720_));
 sky130_fd_sc_hd__o21a_1 _08316_ (.A1(\top.cb_syn.char_path_n[46] ),
    .A2(net202),
    .B1(_04720_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01665_));
 sky130_fd_sc_hd__a221o_1 _08317_ (.A1(\top.cb_syn.char_path_n[46] ),
    .A2(net379),
    .B1(net338),
    .B2(\top.cb_syn.char_path_n[44] ),
    .C1(net182),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04721_));
 sky130_fd_sc_hd__o21a_1 _08318_ (.A1(\top.cb_syn.char_path_n[45] ),
    .A2(net200),
    .B1(_04721_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01664_));
 sky130_fd_sc_hd__a221o_1 _08319_ (.A1(\top.cb_syn.char_path_n[45] ),
    .A2(net381),
    .B1(net338),
    .B2(\top.cb_syn.char_path_n[43] ),
    .C1(net184),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04722_));
 sky130_fd_sc_hd__o21a_1 _08320_ (.A1(\top.cb_syn.char_path_n[44] ),
    .A2(net202),
    .B1(_04722_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01663_));
 sky130_fd_sc_hd__a221o_1 _08321_ (.A1(\top.cb_syn.char_path_n[44] ),
    .A2(net381),
    .B1(net338),
    .B2(\top.cb_syn.char_path_n[42] ),
    .C1(net184),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04723_));
 sky130_fd_sc_hd__o21a_1 _08322_ (.A1(\top.cb_syn.char_path_n[43] ),
    .A2(net202),
    .B1(_04723_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01662_));
 sky130_fd_sc_hd__a221o_1 _08323_ (.A1(\top.cb_syn.char_path_n[43] ),
    .A2(net381),
    .B1(net338),
    .B2(\top.cb_syn.char_path_n[41] ),
    .C1(net184),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04724_));
 sky130_fd_sc_hd__o21a_1 _08324_ (.A1(net1716),
    .A2(net202),
    .B1(_04724_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01661_));
 sky130_fd_sc_hd__a221o_1 _08325_ (.A1(\top.cb_syn.char_path_n[42] ),
    .A2(net379),
    .B1(net336),
    .B2(\top.cb_syn.char_path_n[40] ),
    .C1(net182),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04725_));
 sky130_fd_sc_hd__o21a_1 _08326_ (.A1(\top.cb_syn.char_path_n[41] ),
    .A2(net200),
    .B1(_04725_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01660_));
 sky130_fd_sc_hd__a221o_1 _08327_ (.A1(\top.cb_syn.char_path_n[41] ),
    .A2(net379),
    .B1(net336),
    .B2(\top.cb_syn.char_path_n[39] ),
    .C1(net182),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04726_));
 sky130_fd_sc_hd__o21a_1 _08328_ (.A1(\top.cb_syn.char_path_n[40] ),
    .A2(net200),
    .B1(_04726_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01659_));
 sky130_fd_sc_hd__a221o_1 _08329_ (.A1(\top.cb_syn.char_path_n[40] ),
    .A2(net380),
    .B1(net337),
    .B2(\top.cb_syn.char_path_n[38] ),
    .C1(net183),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04727_));
 sky130_fd_sc_hd__o21a_1 _08330_ (.A1(\top.cb_syn.char_path_n[39] ),
    .A2(net201),
    .B1(_04727_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01658_));
 sky130_fd_sc_hd__a221o_1 _08331_ (.A1(\top.cb_syn.char_path_n[39] ),
    .A2(net380),
    .B1(net337),
    .B2(\top.cb_syn.char_path_n[37] ),
    .C1(net183),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04728_));
 sky130_fd_sc_hd__o21a_1 _08332_ (.A1(\top.cb_syn.char_path_n[38] ),
    .A2(net201),
    .B1(_04728_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01657_));
 sky130_fd_sc_hd__a221o_1 _08333_ (.A1(\top.cb_syn.char_path_n[38] ),
    .A2(net379),
    .B1(net336),
    .B2(\top.cb_syn.char_path_n[36] ),
    .C1(net182),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04729_));
 sky130_fd_sc_hd__o21a_1 _08334_ (.A1(\top.cb_syn.char_path_n[37] ),
    .A2(net200),
    .B1(_04729_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01656_));
 sky130_fd_sc_hd__a221o_1 _08335_ (.A1(\top.cb_syn.char_path_n[37] ),
    .A2(net379),
    .B1(net336),
    .B2(\top.cb_syn.char_path_n[35] ),
    .C1(net182),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04730_));
 sky130_fd_sc_hd__o21a_1 _08336_ (.A1(\top.cb_syn.char_path_n[36] ),
    .A2(net200),
    .B1(_04730_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01655_));
 sky130_fd_sc_hd__a221o_1 _08337_ (.A1(\top.cb_syn.char_path_n[36] ),
    .A2(net379),
    .B1(net336),
    .B2(\top.cb_syn.char_path_n[34] ),
    .C1(net182),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04731_));
 sky130_fd_sc_hd__o21a_1 _08338_ (.A1(\top.cb_syn.char_path_n[35] ),
    .A2(net200),
    .B1(_04731_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01654_));
 sky130_fd_sc_hd__a221o_1 _08339_ (.A1(\top.cb_syn.char_path_n[35] ),
    .A2(net379),
    .B1(net332),
    .B2(\top.cb_syn.char_path_n[33] ),
    .C1(net182),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04732_));
 sky130_fd_sc_hd__o21a_1 _08340_ (.A1(\top.cb_syn.char_path_n[34] ),
    .A2(net200),
    .B1(_04732_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01653_));
 sky130_fd_sc_hd__a221o_1 _08341_ (.A1(\top.cb_syn.char_path_n[34] ),
    .A2(net372),
    .B1(net329),
    .B2(\top.cb_syn.char_path_n[32] ),
    .C1(net177),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04733_));
 sky130_fd_sc_hd__o21a_1 _08342_ (.A1(\top.cb_syn.char_path_n[33] ),
    .A2(net195),
    .B1(_04733_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01652_));
 sky130_fd_sc_hd__a221o_1 _08343_ (.A1(\top.cb_syn.char_path_n[33] ),
    .A2(net371),
    .B1(net328),
    .B2(\top.cb_syn.char_path_n[31] ),
    .C1(net175),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04734_));
 sky130_fd_sc_hd__o21a_1 _08344_ (.A1(\top.cb_syn.char_path_n[32] ),
    .A2(net193),
    .B1(_04734_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01651_));
 sky130_fd_sc_hd__a221o_1 _08345_ (.A1(\top.cb_syn.char_path_n[32] ),
    .A2(net373),
    .B1(net327),
    .B2(\top.cb_syn.char_path_n[30] ),
    .C1(net176),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04735_));
 sky130_fd_sc_hd__o21a_1 _08346_ (.A1(\top.cb_syn.char_path_n[31] ),
    .A2(net194),
    .B1(_04735_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01650_));
 sky130_fd_sc_hd__a221o_1 _08347_ (.A1(\top.cb_syn.char_path_n[31] ),
    .A2(net369),
    .B1(net327),
    .B2(\top.cb_syn.char_path_n[29] ),
    .C1(net173),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04736_));
 sky130_fd_sc_hd__o21a_1 _08348_ (.A1(\top.cb_syn.char_path_n[30] ),
    .A2(net191),
    .B1(_04736_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01649_));
 sky130_fd_sc_hd__a221o_1 _08349_ (.A1(\top.cb_syn.char_path_n[30] ),
    .A2(net373),
    .B1(net327),
    .B2(\top.cb_syn.char_path_n[28] ),
    .C1(net172),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04737_));
 sky130_fd_sc_hd__o21a_1 _08350_ (.A1(net1754),
    .A2(net194),
    .B1(_04737_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01648_));
 sky130_fd_sc_hd__a221o_1 _08351_ (.A1(\top.cb_syn.char_path_n[29] ),
    .A2(net369),
    .B1(net327),
    .B2(\top.cb_syn.char_path_n[27] ),
    .C1(net173),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04738_));
 sky130_fd_sc_hd__o21a_1 _08352_ (.A1(\top.cb_syn.char_path_n[28] ),
    .A2(net190),
    .B1(_04738_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01647_));
 sky130_fd_sc_hd__a221o_1 _08353_ (.A1(\top.cb_syn.char_path_n[28] ),
    .A2(net373),
    .B1(net327),
    .B2(\top.cb_syn.char_path_n[26] ),
    .C1(net176),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04739_));
 sky130_fd_sc_hd__o21a_1 _08354_ (.A1(\top.cb_syn.char_path_n[27] ),
    .A2(net194),
    .B1(_04739_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01646_));
 sky130_fd_sc_hd__a221o_1 _08355_ (.A1(\top.cb_syn.char_path_n[27] ),
    .A2(net373),
    .B1(net327),
    .B2(\top.cb_syn.char_path_n[25] ),
    .C1(net176),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04740_));
 sky130_fd_sc_hd__o21a_1 _08356_ (.A1(\top.cb_syn.char_path_n[26] ),
    .A2(net194),
    .B1(_04740_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01645_));
 sky130_fd_sc_hd__a221o_1 _08357_ (.A1(\top.cb_syn.char_path_n[26] ),
    .A2(net374),
    .B1(net330),
    .B2(\top.cb_syn.char_path_n[24] ),
    .C1(net176),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04741_));
 sky130_fd_sc_hd__o21a_1 _08358_ (.A1(net1781),
    .A2(net194),
    .B1(_04741_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01644_));
 sky130_fd_sc_hd__a221o_1 _08359_ (.A1(\top.cb_syn.char_path_n[25] ),
    .A2(net374),
    .B1(net330),
    .B2(\top.cb_syn.char_path_n[23] ),
    .C1(net177),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04742_));
 sky130_fd_sc_hd__o21a_1 _08360_ (.A1(\top.cb_syn.char_path_n[24] ),
    .A2(net195),
    .B1(_04742_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01643_));
 sky130_fd_sc_hd__a221o_1 _08361_ (.A1(\top.cb_syn.char_path_n[24] ),
    .A2(net373),
    .B1(net330),
    .B2(\top.cb_syn.char_path_n[22] ),
    .C1(net176),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04743_));
 sky130_fd_sc_hd__o21a_1 _08362_ (.A1(\top.cb_syn.char_path_n[23] ),
    .A2(net195),
    .B1(_04743_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01642_));
 sky130_fd_sc_hd__a221o_1 _08363_ (.A1(\top.cb_syn.char_path_n[23] ),
    .A2(net373),
    .B1(net330),
    .B2(\top.cb_syn.char_path_n[21] ),
    .C1(net176),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04744_));
 sky130_fd_sc_hd__o21a_1 _08364_ (.A1(net1766),
    .A2(net195),
    .B1(_04744_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01641_));
 sky130_fd_sc_hd__a221o_1 _08365_ (.A1(\top.cb_syn.char_path_n[22] ),
    .A2(net377),
    .B1(net330),
    .B2(\top.cb_syn.char_path_n[20] ),
    .C1(net177),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04745_));
 sky130_fd_sc_hd__o21a_1 _08366_ (.A1(\top.cb_syn.char_path_n[21] ),
    .A2(net194),
    .B1(_04745_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01640_));
 sky130_fd_sc_hd__a221o_1 _08367_ (.A1(\top.cb_syn.char_path_n[21] ),
    .A2(net377),
    .B1(net330),
    .B2(\top.cb_syn.char_path_n[19] ),
    .C1(net180),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04746_));
 sky130_fd_sc_hd__o21a_1 _08368_ (.A1(\top.cb_syn.char_path_n[20] ),
    .A2(net198),
    .B1(_04746_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01639_));
 sky130_fd_sc_hd__a221o_1 _08369_ (.A1(\top.cb_syn.char_path_n[20] ),
    .A2(net377),
    .B1(net334),
    .B2(\top.cb_syn.char_path_n[18] ),
    .C1(net180),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04747_));
 sky130_fd_sc_hd__o21a_1 _08370_ (.A1(\top.cb_syn.char_path_n[19] ),
    .A2(net198),
    .B1(_04747_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01638_));
 sky130_fd_sc_hd__a221o_1 _08371_ (.A1(\top.cb_syn.char_path_n[19] ),
    .A2(net378),
    .B1(net334),
    .B2(\top.cb_syn.char_path_n[17] ),
    .C1(net181),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04748_));
 sky130_fd_sc_hd__o21a_1 _08372_ (.A1(\top.cb_syn.char_path_n[18] ),
    .A2(net199),
    .B1(_04748_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01637_));
 sky130_fd_sc_hd__a221o_1 _08373_ (.A1(\top.cb_syn.char_path_n[18] ),
    .A2(net378),
    .B1(net335),
    .B2(\top.cb_syn.char_path_n[16] ),
    .C1(net181),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04749_));
 sky130_fd_sc_hd__o21a_1 _08374_ (.A1(net1751),
    .A2(net199),
    .B1(_04749_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01636_));
 sky130_fd_sc_hd__a221o_1 _08375_ (.A1(\top.cb_syn.char_path_n[17] ),
    .A2(net385),
    .B1(net340),
    .B2(\top.cb_syn.char_path_n[15] ),
    .C1(net188),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04750_));
 sky130_fd_sc_hd__o21a_1 _08376_ (.A1(\top.cb_syn.char_path_n[16] ),
    .A2(net205),
    .B1(_04750_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01635_));
 sky130_fd_sc_hd__a221o_1 _08377_ (.A1(\top.cb_syn.char_path_n[16] ),
    .A2(net385),
    .B1(net340),
    .B2(\top.cb_syn.char_path_n[14] ),
    .C1(net188),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04751_));
 sky130_fd_sc_hd__o21a_1 _08378_ (.A1(\top.cb_syn.char_path_n[15] ),
    .A2(net205),
    .B1(_04751_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01634_));
 sky130_fd_sc_hd__a221o_1 _08379_ (.A1(\top.cb_syn.char_path_n[15] ),
    .A2(net384),
    .B1(net340),
    .B2(\top.cb_syn.char_path_n[13] ),
    .C1(net187),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04752_));
 sky130_fd_sc_hd__o21a_1 _08380_ (.A1(\top.cb_syn.char_path_n[14] ),
    .A2(net204),
    .B1(_04752_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01633_));
 sky130_fd_sc_hd__a221o_1 _08381_ (.A1(\top.cb_syn.char_path_n[14] ),
    .A2(net384),
    .B1(net340),
    .B2(\top.cb_syn.char_path_n[12] ),
    .C1(net187),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04753_));
 sky130_fd_sc_hd__o21a_1 _08382_ (.A1(\top.cb_syn.char_path_n[13] ),
    .A2(net204),
    .B1(_04753_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01632_));
 sky130_fd_sc_hd__a221o_1 _08383_ (.A1(\top.cb_syn.char_path_n[13] ),
    .A2(net383),
    .B1(net340),
    .B2(\top.cb_syn.char_path_n[11] ),
    .C1(net187),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04754_));
 sky130_fd_sc_hd__o21a_1 _08384_ (.A1(\top.cb_syn.char_path_n[12] ),
    .A2(net204),
    .B1(_04754_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01631_));
 sky130_fd_sc_hd__a221o_1 _08385_ (.A1(\top.cb_syn.char_path_n[12] ),
    .A2(net383),
    .B1(net340),
    .B2(\top.cb_syn.char_path_n[10] ),
    .C1(net187),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04755_));
 sky130_fd_sc_hd__o21a_1 _08386_ (.A1(net1782),
    .A2(net204),
    .B1(_04755_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01630_));
 sky130_fd_sc_hd__a221o_1 _08387_ (.A1(\top.cb_syn.char_path_n[11] ),
    .A2(net383),
    .B1(net339),
    .B2(\top.cb_syn.char_path_n[9] ),
    .C1(net186),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04756_));
 sky130_fd_sc_hd__o21a_1 _08388_ (.A1(\top.cb_syn.char_path_n[10] ),
    .A2(net203),
    .B1(_04756_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01629_));
 sky130_fd_sc_hd__a221o_1 _08389_ (.A1(\top.cb_syn.char_path_n[10] ),
    .A2(net380),
    .B1(net337),
    .B2(\top.cb_syn.char_path_n[8] ),
    .C1(net183),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04757_));
 sky130_fd_sc_hd__o21a_1 _08390_ (.A1(\top.cb_syn.char_path_n[9] ),
    .A2(net202),
    .B1(_04757_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01628_));
 sky130_fd_sc_hd__a221o_1 _08391_ (.A1(\top.cb_syn.char_path_n[9] ),
    .A2(net381),
    .B1(net337),
    .B2(\top.cb_syn.char_path_n[7] ),
    .C1(net184),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04758_));
 sky130_fd_sc_hd__o21a_1 _08392_ (.A1(\top.cb_syn.char_path_n[8] ),
    .A2(net201),
    .B1(_04758_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01627_));
 sky130_fd_sc_hd__a221o_1 _08393_ (.A1(\top.cb_syn.char_path_n[8] ),
    .A2(net376),
    .B1(net333),
    .B2(\top.cb_syn.char_path_n[6] ),
    .C1(net179),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04759_));
 sky130_fd_sc_hd__o21a_1 _08394_ (.A1(\top.cb_syn.char_path_n[7] ),
    .A2(net197),
    .B1(_04759_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01626_));
 sky130_fd_sc_hd__a221o_1 _08395_ (.A1(\top.cb_syn.char_path_n[7] ),
    .A2(net375),
    .B1(net332),
    .B2(\top.cb_syn.char_path_n[5] ),
    .C1(net178),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04760_));
 sky130_fd_sc_hd__o21a_1 _08396_ (.A1(\top.cb_syn.char_path_n[6] ),
    .A2(net196),
    .B1(_04760_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01625_));
 sky130_fd_sc_hd__a221o_1 _08397_ (.A1(\top.cb_syn.char_path_n[6] ),
    .A2(net375),
    .B1(net332),
    .B2(\top.cb_syn.char_path_n[4] ),
    .C1(net178),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04761_));
 sky130_fd_sc_hd__o21a_1 _08398_ (.A1(\top.cb_syn.char_path_n[5] ),
    .A2(net197),
    .B1(_04761_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01624_));
 sky130_fd_sc_hd__a221o_1 _08399_ (.A1(\top.cb_syn.char_path_n[5] ),
    .A2(net375),
    .B1(net332),
    .B2(\top.cb_syn.char_path_n[3] ),
    .C1(net178),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04762_));
 sky130_fd_sc_hd__o21a_1 _08400_ (.A1(\top.cb_syn.char_path_n[4] ),
    .A2(net196),
    .B1(_04762_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01623_));
 sky130_fd_sc_hd__a221o_1 _08401_ (.A1(\top.cb_syn.char_path_n[4] ),
    .A2(net375),
    .B1(net332),
    .B2(\top.cb_syn.char_path_n[2] ),
    .C1(net179),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04763_));
 sky130_fd_sc_hd__o21a_1 _08402_ (.A1(\top.cb_syn.char_path_n[3] ),
    .A2(net197),
    .B1(_04763_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01622_));
 sky130_fd_sc_hd__a221o_1 _08403_ (.A1(\top.cb_syn.char_path_n[3] ),
    .A2(net376),
    .B1(net332),
    .B2(\top.cb_syn.char_path_n[1] ),
    .C1(net179),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04764_));
 sky130_fd_sc_hd__o21a_1 _08404_ (.A1(\top.cb_syn.char_path_n[2] ),
    .A2(net197),
    .B1(_04764_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01621_));
 sky130_fd_sc_hd__a211o_1 _08405_ (.A1(\top.cb_syn.char_path_n[2] ),
    .A2(net370),
    .B1(net174),
    .C1(net520),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04765_));
 sky130_fd_sc_hd__o21a_1 _08406_ (.A1(\top.cb_syn.char_path_n[1] ),
    .A2(net192),
    .B1(_04765_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01620_));
 sky130_fd_sc_hd__o211a_1 _08407_ (.A1(net522),
    .A2(net523),
    .B1(_04559_),
    .C1(_04561_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04766_));
 sky130_fd_sc_hd__mux2_1 _08408_ (.A0(net1515),
    .A1(_02554_),
    .S(_04766_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01619_));
 sky130_fd_sc_hd__nor2_1 _08409_ (.A(_02885_),
    .B(_04606_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04767_));
 sky130_fd_sc_hd__a21o_1 _08410_ (.A1(net488),
    .A2(net519),
    .B1(net424),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04768_));
 sky130_fd_sc_hd__o21bai_2 _08411_ (.A1(net519),
    .A2(net524),
    .B1_N(_04583_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04769_));
 sky130_fd_sc_hd__nor2_1 _08412_ (.A(_04767_),
    .B(_04768_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04770_));
 sky130_fd_sc_hd__or2_1 _08413_ (.A(_04767_),
    .B(_04768_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04771_));
 sky130_fd_sc_hd__nor2_4 _08414_ (.A(_04769_),
    .B(_04771_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04772_));
 sky130_fd_sc_hd__mux2_1 _08415_ (.A0(\top.cb_syn.h_element[62] ),
    .A1(\top.cb_syn.h_element[53] ),
    .S(net518),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04773_));
 sky130_fd_sc_hd__mux2_1 _08416_ (.A0(net1050),
    .A1(_04773_),
    .S(_04772_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01618_));
 sky130_fd_sc_hd__mux2_1 _08417_ (.A0(\top.cb_syn.h_element[61] ),
    .A1(\top.cb_syn.h_element[52] ),
    .S(net517),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04774_));
 sky130_fd_sc_hd__mux2_1 _08418_ (.A0(\top.cb_syn.char_index[6] ),
    .A1(_04774_),
    .S(_04772_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01617_));
 sky130_fd_sc_hd__mux2_1 _08419_ (.A0(\top.cb_syn.h_element[60] ),
    .A1(\top.cb_syn.h_element[51] ),
    .S(net518),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04775_));
 sky130_fd_sc_hd__mux2_1 _08420_ (.A0(\top.cb_syn.char_index[5] ),
    .A1(_04775_),
    .S(_04772_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01616_));
 sky130_fd_sc_hd__mux2_1 _08421_ (.A0(\top.cb_syn.h_element[59] ),
    .A1(\top.cb_syn.h_element[50] ),
    .S(net517),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04776_));
 sky130_fd_sc_hd__mux2_1 _08422_ (.A0(\top.cb_syn.char_index[4] ),
    .A1(_04776_),
    .S(_04772_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01615_));
 sky130_fd_sc_hd__mux2_1 _08423_ (.A0(\top.cb_syn.h_element[58] ),
    .A1(\top.cb_syn.h_element[49] ),
    .S(net517),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04777_));
 sky130_fd_sc_hd__mux2_1 _08424_ (.A0(\top.cb_syn.char_index[3] ),
    .A1(_04777_),
    .S(_04772_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01614_));
 sky130_fd_sc_hd__mux2_1 _08425_ (.A0(\top.cb_syn.h_element[57] ),
    .A1(\top.cb_syn.h_element[48] ),
    .S(net517),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04778_));
 sky130_fd_sc_hd__mux2_1 _08426_ (.A0(\top.cb_syn.char_index[2] ),
    .A1(_04778_),
    .S(_04772_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01613_));
 sky130_fd_sc_hd__mux2_1 _08427_ (.A0(\top.cb_syn.h_element[56] ),
    .A1(\top.cb_syn.h_element[47] ),
    .S(net517),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04779_));
 sky130_fd_sc_hd__mux2_1 _08428_ (.A0(\top.cb_syn.char_index[1] ),
    .A1(_04779_),
    .S(_04772_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01612_));
 sky130_fd_sc_hd__mux2_1 _08429_ (.A0(\top.cb_syn.h_element[55] ),
    .A1(\top.cb_syn.h_element[46] ),
    .S(net517),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04780_));
 sky130_fd_sc_hd__mux2_1 _08430_ (.A0(\top.cb_syn.char_index[0] ),
    .A1(_04780_),
    .S(_04772_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01611_));
 sky130_fd_sc_hd__nor3b_1 _08431_ (.A(_04586_),
    .B(_04610_),
    .C_N(_04178_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04781_));
 sky130_fd_sc_hd__mux2_1 _08432_ (.A0(net1119),
    .A1(\top.cb_syn.char_path_n[127] ),
    .S(net230),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01610_));
 sky130_fd_sc_hd__mux2_1 _08433_ (.A0(net1139),
    .A1(\top.cb_syn.char_path_n[126] ),
    .S(net230),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01609_));
 sky130_fd_sc_hd__mux2_1 _08434_ (.A0(net1413),
    .A1(\top.cb_syn.char_path_n[125] ),
    .S(net230),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01608_));
 sky130_fd_sc_hd__mux2_1 _08435_ (.A0(net1303),
    .A1(\top.cb_syn.char_path_n[124] ),
    .S(net230),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01607_));
 sky130_fd_sc_hd__mux2_1 _08436_ (.A0(net1333),
    .A1(\top.cb_syn.char_path_n[123] ),
    .S(net234),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01606_));
 sky130_fd_sc_hd__mux2_1 _08437_ (.A0(net1280),
    .A1(\top.cb_syn.char_path_n[122] ),
    .S(net234),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01605_));
 sky130_fd_sc_hd__mux2_1 _08438_ (.A0(net1317),
    .A1(\top.cb_syn.char_path_n[121] ),
    .S(net234),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01604_));
 sky130_fd_sc_hd__mux2_1 _08439_ (.A0(net1079),
    .A1(\top.cb_syn.char_path_n[120] ),
    .S(net235),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01603_));
 sky130_fd_sc_hd__mux2_1 _08440_ (.A0(net1099),
    .A1(\top.cb_syn.char_path_n[119] ),
    .S(net235),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01602_));
 sky130_fd_sc_hd__mux2_1 _08441_ (.A0(net1088),
    .A1(\top.cb_syn.char_path_n[118] ),
    .S(net235),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01601_));
 sky130_fd_sc_hd__mux2_1 _08442_ (.A0(net1272),
    .A1(\top.cb_syn.char_path_n[117] ),
    .S(net235),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01600_));
 sky130_fd_sc_hd__mux2_1 _08443_ (.A0(net1161),
    .A1(\top.cb_syn.char_path_n[116] ),
    .S(net242),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01599_));
 sky130_fd_sc_hd__mux2_1 _08444_ (.A0(net1133),
    .A1(\top.cb_syn.char_path_n[115] ),
    .S(net242),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01598_));
 sky130_fd_sc_hd__mux2_1 _08445_ (.A0(net1277),
    .A1(\top.cb_syn.char_path_n[114] ),
    .S(net242),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01597_));
 sky130_fd_sc_hd__mux2_1 _08446_ (.A0(net1149),
    .A1(\top.cb_syn.char_path_n[113] ),
    .S(net243),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01596_));
 sky130_fd_sc_hd__mux2_1 _08447_ (.A0(net1061),
    .A1(\top.cb_syn.char_path_n[112] ),
    .S(net242),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01595_));
 sky130_fd_sc_hd__mux2_1 _08448_ (.A0(net1097),
    .A1(\top.cb_syn.char_path_n[111] ),
    .S(net242),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01594_));
 sky130_fd_sc_hd__mux2_1 _08449_ (.A0(net1063),
    .A1(\top.cb_syn.char_path_n[110] ),
    .S(net244),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01593_));
 sky130_fd_sc_hd__mux2_1 _08450_ (.A0(net1266),
    .A1(\top.cb_syn.char_path_n[109] ),
    .S(net244),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01592_));
 sky130_fd_sc_hd__mux2_1 _08451_ (.A0(net1210),
    .A1(\top.cb_syn.char_path_n[108] ),
    .S(net244),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01591_));
 sky130_fd_sc_hd__mux2_1 _08452_ (.A0(net1370),
    .A1(\top.cb_syn.char_path_n[107] ),
    .S(net244),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01590_));
 sky130_fd_sc_hd__mux2_1 _08453_ (.A0(net1358),
    .A1(\top.cb_syn.char_path_n[106] ),
    .S(net241),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01589_));
 sky130_fd_sc_hd__mux2_1 _08454_ (.A0(net1115),
    .A1(\top.cb_syn.char_path_n[105] ),
    .S(net240),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01588_));
 sky130_fd_sc_hd__mux2_1 _08455_ (.A0(net1238),
    .A1(\top.cb_syn.char_path_n[104] ),
    .S(net240),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01587_));
 sky130_fd_sc_hd__mux2_1 _08456_ (.A0(net1203),
    .A1(\top.cb_syn.char_path_n[103] ),
    .S(net239),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01586_));
 sky130_fd_sc_hd__mux2_1 _08457_ (.A0(net1216),
    .A1(\top.cb_syn.char_path_n[102] ),
    .S(net239),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01585_));
 sky130_fd_sc_hd__mux2_1 _08458_ (.A0(net1242),
    .A1(\top.cb_syn.char_path_n[101] ),
    .S(net239),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01584_));
 sky130_fd_sc_hd__mux2_1 _08459_ (.A0(net1213),
    .A1(\top.cb_syn.char_path_n[100] ),
    .S(net239),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01583_));
 sky130_fd_sc_hd__mux2_1 _08460_ (.A0(net1302),
    .A1(\top.cb_syn.char_path_n[99] ),
    .S(net239),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01582_));
 sky130_fd_sc_hd__mux2_1 _08461_ (.A0(net1404),
    .A1(\top.cb_syn.char_path_n[98] ),
    .S(net232),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01581_));
 sky130_fd_sc_hd__mux2_1 _08462_ (.A0(net1320),
    .A1(\top.cb_syn.char_path_n[97] ),
    .S(net237),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01580_));
 sky130_fd_sc_hd__mux2_1 _08463_ (.A0(net1158),
    .A1(\top.cb_syn.char_path_n[96] ),
    .S(net232),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01579_));
 sky130_fd_sc_hd__mux2_1 _08464_ (.A0(net1329),
    .A1(\top.cb_syn.char_path_n[95] ),
    .S(net233),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01578_));
 sky130_fd_sc_hd__mux2_1 _08465_ (.A0(net1074),
    .A1(net1805),
    .S(net230),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01577_));
 sky130_fd_sc_hd__mux2_1 _08466_ (.A0(net1292),
    .A1(\top.cb_syn.char_path_n[93] ),
    .S(net230),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01576_));
 sky130_fd_sc_hd__mux2_1 _08467_ (.A0(net1082),
    .A1(\top.cb_syn.char_path_n[92] ),
    .S(net236),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01575_));
 sky130_fd_sc_hd__mux2_1 _08468_ (.A0(net1439),
    .A1(\top.cb_syn.char_path_n[91] ),
    .S(net236),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01574_));
 sky130_fd_sc_hd__mux2_1 _08469_ (.A0(net1132),
    .A1(\top.cb_syn.char_path_n[90] ),
    .S(net234),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01573_));
 sky130_fd_sc_hd__mux2_1 _08470_ (.A0(net1554),
    .A1(net1808),
    .S(net234),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01572_));
 sky130_fd_sc_hd__mux2_1 _08471_ (.A0(net1186),
    .A1(\top.cb_syn.char_path_n[88] ),
    .S(net236),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01571_));
 sky130_fd_sc_hd__mux2_1 _08472_ (.A0(net1262),
    .A1(\top.cb_syn.char_path_n[87] ),
    .S(net236),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01570_));
 sky130_fd_sc_hd__mux2_1 _08473_ (.A0(net1235),
    .A1(\top.cb_syn.char_path_n[86] ),
    .S(net235),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01569_));
 sky130_fd_sc_hd__mux2_1 _08474_ (.A0(net1269),
    .A1(\top.cb_syn.char_path_n[85] ),
    .S(net235),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01568_));
 sky130_fd_sc_hd__mux2_1 _08475_ (.A0(net1231),
    .A1(\top.cb_syn.char_path_n[84] ),
    .S(net242),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01567_));
 sky130_fd_sc_hd__mux2_1 _08476_ (.A0(net1184),
    .A1(\top.cb_syn.char_path_n[83] ),
    .S(net243),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01566_));
 sky130_fd_sc_hd__mux2_1 _08477_ (.A0(net1264),
    .A1(\top.cb_syn.char_path_n[82] ),
    .S(net246),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01565_));
 sky130_fd_sc_hd__mux2_1 _08478_ (.A0(net1245),
    .A1(\top.cb_syn.char_path_n[81] ),
    .S(net246),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01564_));
 sky130_fd_sc_hd__mux2_1 _08479_ (.A0(net1112),
    .A1(\top.cb_syn.char_path_n[80] ),
    .S(net243),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01563_));
 sky130_fd_sc_hd__mux2_1 _08480_ (.A0(net1197),
    .A1(\top.cb_syn.char_path_n[79] ),
    .S(net243),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01562_));
 sky130_fd_sc_hd__mux2_1 _08481_ (.A0(net1513),
    .A1(\top.cb_syn.char_path_n[78] ),
    .S(net245),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01561_));
 sky130_fd_sc_hd__mux2_1 _08482_ (.A0(net1163),
    .A1(\top.cb_syn.char_path_n[77] ),
    .S(net245),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01560_));
 sky130_fd_sc_hd__mux2_1 _08483_ (.A0(net1539),
    .A1(\top.cb_syn.char_path_n[76] ),
    .S(net245),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01559_));
 sky130_fd_sc_hd__mux2_1 _08484_ (.A0(net1367),
    .A1(\top.cb_syn.char_path_n[75] ),
    .S(net244),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01558_));
 sky130_fd_sc_hd__mux2_1 _08485_ (.A0(net1362),
    .A1(\top.cb_syn.char_path_n[74] ),
    .S(net241),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01557_));
 sky130_fd_sc_hd__mux2_1 _08486_ (.A0(net1176),
    .A1(\top.cb_syn.char_path_n[73] ),
    .S(net240),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01556_));
 sky130_fd_sc_hd__mux2_1 _08487_ (.A0(net1309),
    .A1(\top.cb_syn.char_path_n[72] ),
    .S(net239),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01555_));
 sky130_fd_sc_hd__mux2_1 _08488_ (.A0(net1347),
    .A1(\top.cb_syn.char_path_n[71] ),
    .S(net239),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01554_));
 sky130_fd_sc_hd__mux2_1 _08489_ (.A0(net1177),
    .A1(\top.cb_syn.char_path_n[70] ),
    .S(net237),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01553_));
 sky130_fd_sc_hd__mux2_1 _08490_ (.A0(net1086),
    .A1(\top.cb_syn.char_path_n[69] ),
    .S(net237),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01552_));
 sky130_fd_sc_hd__mux2_1 _08491_ (.A0(net1120),
    .A1(\top.cb_syn.char_path_n[68] ),
    .S(net237),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01551_));
 sky130_fd_sc_hd__mux2_1 _08492_ (.A0(net1094),
    .A1(\top.cb_syn.char_path_n[67] ),
    .S(net237),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01550_));
 sky130_fd_sc_hd__mux2_1 _08493_ (.A0(net1423),
    .A1(\top.cb_syn.char_path_n[66] ),
    .S(net232),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01549_));
 sky130_fd_sc_hd__mux2_1 _08494_ (.A0(net1385),
    .A1(\top.cb_syn.char_path_n[65] ),
    .S(net238),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01548_));
 sky130_fd_sc_hd__mux2_1 _08495_ (.A0(net1225),
    .A1(\top.cb_syn.char_path_n[64] ),
    .S(net230),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01547_));
 sky130_fd_sc_hd__mux2_1 _08496_ (.A0(net1100),
    .A1(\top.cb_syn.char_path_n[63] ),
    .S(net230),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01546_));
 sky130_fd_sc_hd__mux2_1 _08497_ (.A0(net1089),
    .A1(\top.cb_syn.char_path_n[62] ),
    .S(net230),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01545_));
 sky130_fd_sc_hd__mux2_1 _08498_ (.A0(net1295),
    .A1(\top.cb_syn.char_path_n[61] ),
    .S(net230),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01544_));
 sky130_fd_sc_hd__mux2_1 _08499_ (.A0(net1209),
    .A1(\top.cb_syn.char_path_n[60] ),
    .S(net231),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01543_));
 sky130_fd_sc_hd__mux2_1 _08500_ (.A0(net1387),
    .A1(\top.cb_syn.char_path_n[59] ),
    .S(net231),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01542_));
 sky130_fd_sc_hd__mux2_1 _08501_ (.A0(net1291),
    .A1(\top.cb_syn.char_path_n[58] ),
    .S(net231),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01541_));
 sky130_fd_sc_hd__mux2_1 _08502_ (.A0(net1336),
    .A1(\top.cb_syn.char_path_n[57] ),
    .S(net231),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01540_));
 sky130_fd_sc_hd__mux2_1 _08503_ (.A0(net1087),
    .A1(\top.cb_syn.char_path_n[56] ),
    .S(net233),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01539_));
 sky130_fd_sc_hd__mux2_1 _08504_ (.A0(net1151),
    .A1(\top.cb_syn.char_path_n[55] ),
    .S(net232),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01538_));
 sky130_fd_sc_hd__mux2_1 _08505_ (.A0(net1221),
    .A1(\top.cb_syn.char_path_n[54] ),
    .S(net232),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01537_));
 sky130_fd_sc_hd__mux2_1 _08506_ (.A0(net1071),
    .A1(\top.cb_syn.char_path_n[53] ),
    .S(net232),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01536_));
 sky130_fd_sc_hd__mux2_1 _08507_ (.A0(net1136),
    .A1(\top.cb_syn.char_path_n[52] ),
    .S(net242),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01535_));
 sky130_fd_sc_hd__mux2_1 _08508_ (.A0(net1121),
    .A1(\top.cb_syn.char_path_n[51] ),
    .S(net242),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01534_));
 sky130_fd_sc_hd__mux2_1 _08509_ (.A0(net1129),
    .A1(\top.cb_syn.char_path_n[50] ),
    .S(net242),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01533_));
 sky130_fd_sc_hd__mux2_1 _08510_ (.A0(net1416),
    .A1(\top.cb_syn.char_path_n[49] ),
    .S(net243),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01532_));
 sky130_fd_sc_hd__mux2_1 _08511_ (.A0(net1310),
    .A1(\top.cb_syn.char_path_n[48] ),
    .S(net243),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01531_));
 sky130_fd_sc_hd__mux2_1 _08512_ (.A0(net1157),
    .A1(\top.cb_syn.char_path_n[47] ),
    .S(net242),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01530_));
 sky130_fd_sc_hd__mux2_1 _08513_ (.A0(net1067),
    .A1(\top.cb_syn.char_path_n[46] ),
    .S(net244),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01529_));
 sky130_fd_sc_hd__mux2_1 _08514_ (.A0(net1255),
    .A1(\top.cb_syn.char_path_n[45] ),
    .S(net244),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01528_));
 sky130_fd_sc_hd__mux2_1 _08515_ (.A0(net1322),
    .A1(\top.cb_syn.char_path_n[44] ),
    .S(net244),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01527_));
 sky130_fd_sc_hd__mux2_1 _08516_ (.A0(net1402),
    .A1(\top.cb_syn.char_path_n[43] ),
    .S(net244),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01526_));
 sky130_fd_sc_hd__mux2_1 _08517_ (.A0(net1360),
    .A1(\top.cb_syn.char_path_n[42] ),
    .S(net241),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01525_));
 sky130_fd_sc_hd__mux2_1 _08518_ (.A0(net1357),
    .A1(\top.cb_syn.char_path_n[41] ),
    .S(net240),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01524_));
 sky130_fd_sc_hd__mux2_1 _08519_ (.A0(net1319),
    .A1(\top.cb_syn.char_path_n[40] ),
    .S(net240),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01523_));
 sky130_fd_sc_hd__mux2_1 _08520_ (.A0(net1349),
    .A1(\top.cb_syn.char_path_n[39] ),
    .S(net239),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01522_));
 sky130_fd_sc_hd__mux2_1 _08521_ (.A0(net1298),
    .A1(\top.cb_syn.char_path_n[38] ),
    .S(net239),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01521_));
 sky130_fd_sc_hd__mux2_1 _08522_ (.A0(net1271),
    .A1(\top.cb_syn.char_path_n[37] ),
    .S(net239),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01520_));
 sky130_fd_sc_hd__mux2_1 _08523_ (.A0(net1141),
    .A1(\top.cb_syn.char_path_n[36] ),
    .S(net237),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01519_));
 sky130_fd_sc_hd__mux2_1 _08524_ (.A0(net1111),
    .A1(\top.cb_syn.char_path_n[35] ),
    .S(net238),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01518_));
 sky130_fd_sc_hd__mux2_1 _08525_ (.A0(net1354),
    .A1(\top.cb_syn.char_path_n[34] ),
    .S(net232),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01517_));
 sky130_fd_sc_hd__mux2_1 _08526_ (.A0(net1324),
    .A1(\top.cb_syn.char_path_n[33] ),
    .S(net237),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01516_));
 sky130_fd_sc_hd__mux2_1 _08527_ (.A0(net1193),
    .A1(\top.cb_syn.char_path_n[32] ),
    .S(net232),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01515_));
 sky130_fd_sc_hd__mux2_1 _08528_ (.A0(net1297),
    .A1(\top.cb_syn.char_path_n[31] ),
    .S(net231),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01514_));
 sky130_fd_sc_hd__mux2_1 _08529_ (.A0(net1152),
    .A1(\top.cb_syn.char_path_n[30] ),
    .S(net234),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01513_));
 sky130_fd_sc_hd__mux2_1 _08530_ (.A0(net1426),
    .A1(\top.cb_syn.char_path_n[29] ),
    .S(net234),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01512_));
 sky130_fd_sc_hd__mux2_1 _08531_ (.A0(net1068),
    .A1(\top.cb_syn.char_path_n[28] ),
    .S(net234),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01511_));
 sky130_fd_sc_hd__mux2_1 _08532_ (.A0(net1384),
    .A1(\top.cb_syn.char_path_n[27] ),
    .S(net234),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01510_));
 sky130_fd_sc_hd__mux2_1 _08533_ (.A0(net1128),
    .A1(\top.cb_syn.char_path_n[26] ),
    .S(net236),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01509_));
 sky130_fd_sc_hd__mux2_1 _08534_ (.A0(net1342),
    .A1(\top.cb_syn.char_path_n[25] ),
    .S(net234),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01508_));
 sky130_fd_sc_hd__mux2_1 _08535_ (.A0(net1230),
    .A1(\top.cb_syn.char_path_n[24] ),
    .S(net235),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01507_));
 sky130_fd_sc_hd__mux2_1 _08536_ (.A0(net1056),
    .A1(\top.cb_syn.char_path_n[23] ),
    .S(net236),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01506_));
 sky130_fd_sc_hd__mux2_1 _08537_ (.A0(net1304),
    .A1(\top.cb_syn.char_path_n[22] ),
    .S(net235),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01505_));
 sky130_fd_sc_hd__mux2_1 _08538_ (.A0(net1171),
    .A1(\top.cb_syn.char_path_n[21] ),
    .S(net235),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01504_));
 sky130_fd_sc_hd__mux2_1 _08539_ (.A0(net1220),
    .A1(\top.cb_syn.char_path_n[20] ),
    .S(net235),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01503_));
 sky130_fd_sc_hd__mux2_1 _08540_ (.A0(net1228),
    .A1(\top.cb_syn.char_path_n[19] ),
    .S(net246),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01502_));
 sky130_fd_sc_hd__mux2_1 _08541_ (.A0(net1170),
    .A1(\top.cb_syn.char_path_n[18] ),
    .S(net246),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01501_));
 sky130_fd_sc_hd__mux2_1 _08542_ (.A0(net1198),
    .A1(\top.cb_syn.char_path_n[17] ),
    .S(net243),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01500_));
 sky130_fd_sc_hd__mux2_1 _08543_ (.A0(net1104),
    .A1(\top.cb_syn.char_path_n[16] ),
    .S(net243),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01499_));
 sky130_fd_sc_hd__mux2_1 _08544_ (.A0(net1080),
    .A1(\top.cb_syn.char_path_n[15] ),
    .S(net243),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01498_));
 sky130_fd_sc_hd__mux2_1 _08545_ (.A0(net1179),
    .A1(\top.cb_syn.char_path_n[14] ),
    .S(net245),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01497_));
 sky130_fd_sc_hd__mux2_1 _08546_ (.A0(net1123),
    .A1(\top.cb_syn.char_path_n[13] ),
    .S(net245),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01496_));
 sky130_fd_sc_hd__mux2_1 _08547_ (.A0(net1287),
    .A1(\top.cb_syn.char_path_n[12] ),
    .S(net245),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01495_));
 sky130_fd_sc_hd__mux2_1 _08548_ (.A0(net1241),
    .A1(\top.cb_syn.char_path_n[11] ),
    .S(net244),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01494_));
 sky130_fd_sc_hd__mux2_1 _08549_ (.A0(net1321),
    .A1(\top.cb_syn.char_path_n[10] ),
    .S(net240),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01493_));
 sky130_fd_sc_hd__mux2_1 _08550_ (.A0(net1368),
    .A1(\top.cb_syn.char_path_n[9] ),
    .S(net240),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01492_));
 sky130_fd_sc_hd__mux2_1 _08551_ (.A0(net1323),
    .A1(\top.cb_syn.char_path_n[8] ),
    .S(net240),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01491_));
 sky130_fd_sc_hd__mux2_1 _08552_ (.A0(net1284),
    .A1(\top.cb_syn.char_path_n[7] ),
    .S(net240),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01490_));
 sky130_fd_sc_hd__mux2_1 _08553_ (.A0(net1327),
    .A1(\top.cb_syn.char_path_n[6] ),
    .S(net238),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01489_));
 sky130_fd_sc_hd__mux2_1 _08554_ (.A0(net1420),
    .A1(\top.cb_syn.char_path_n[5] ),
    .S(net237),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01488_));
 sky130_fd_sc_hd__mux2_1 _08555_ (.A0(net1334),
    .A1(\top.cb_syn.char_path_n[4] ),
    .S(net237),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01487_));
 sky130_fd_sc_hd__mux2_1 _08556_ (.A0(net1182),
    .A1(\top.cb_syn.char_path_n[3] ),
    .S(net237),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01486_));
 sky130_fd_sc_hd__mux2_1 _08557_ (.A0(net1409),
    .A1(\top.cb_syn.char_path_n[2] ),
    .S(net232),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01485_));
 sky130_fd_sc_hd__mux2_1 _08558_ (.A0(net1090),
    .A1(\top.cb_syn.char_path_n[1] ),
    .S(net238),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01484_));
 sky130_fd_sc_hd__mux2_1 _08559_ (.A0(net1153),
    .A1(\top.cb_syn.char_path_n[0] ),
    .S(net232),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01483_));
 sky130_fd_sc_hd__o311a_1 _08560_ (.A1(net515),
    .A2(\top.cb_syn.curr_state[5] ),
    .A3(_04178_),
    .B1(_04607_),
    .C1(net464),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04782_));
 sky130_fd_sc_hd__or3b_1 _08561_ (.A(_04197_),
    .B(_04609_),
    .C_N(_04782_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04783_));
 sky130_fd_sc_hd__or4_1 _08562_ (.A(net519),
    .B(net515),
    .C(\top.cb_syn.curr_state[5] ),
    .D(_02895_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04784_));
 sky130_fd_sc_hd__nand2_1 _08563_ (.A(_04195_),
    .B(_04784_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04785_));
 sky130_fd_sc_hd__mux2_1 _08564_ (.A0(_04785_),
    .A1(net491),
    .S(_04783_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01482_));
 sky130_fd_sc_hd__or3_1 _08565_ (.A(_02543_),
    .B(\top.cb_syn.h_element[63] ),
    .C(_04562_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04786_));
 sky130_fd_sc_hd__o21a_1 _08566_ (.A1(_02538_),
    .A2(net515),
    .B1(_04786_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04787_));
 sky130_fd_sc_hd__or3_1 _08567_ (.A(_04202_),
    .B(_04771_),
    .C(_04787_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04788_));
 sky130_fd_sc_hd__mux2_1 _08568_ (.A0(_02538_),
    .A1(net1541),
    .S(_04788_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01481_));
 sky130_fd_sc_hd__nor2_1 _08569_ (.A(net496),
    .B(net498),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04789_));
 sky130_fd_sc_hd__or4_1 _08570_ (.A(\top.cb_syn.end_cnt[3] ),
    .B(net493),
    .C(net496),
    .D(net498),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04790_));
 sky130_fd_sc_hd__or3_2 _08571_ (.A(\top.cb_syn.end_cnt[5] ),
    .B(\top.cb_syn.end_cnt[4] ),
    .C(_04790_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04791_));
 sky130_fd_sc_hd__o22ai_2 _08572_ (.A1(_04199_),
    .A2(_04630_),
    .B1(_04791_),
    .B2(\top.cb_syn.end_cnt[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04792_));
 sky130_fd_sc_hd__mux4_1 _08573_ (.A0(\top.cb_syn.char_path_n[81] ),
    .A1(\top.cb_syn.char_path_n[82] ),
    .A2(\top.cb_syn.char_path_n[85] ),
    .A3(\top.cb_syn.char_path_n[86] ),
    .S0(net501),
    .S1(net495),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04793_));
 sky130_fd_sc_hd__mux4_1 _08574_ (.A0(\top.cb_syn.char_path_n[83] ),
    .A1(\top.cb_syn.char_path_n[84] ),
    .A2(\top.cb_syn.char_path_n[87] ),
    .A3(\top.cb_syn.char_path_n[88] ),
    .S0(net501),
    .S1(net495),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04794_));
 sky130_fd_sc_hd__mux2_1 _08575_ (.A0(_04793_),
    .A1(_04794_),
    .S(net496),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04795_));
 sky130_fd_sc_hd__mux4_1 _08576_ (.A0(\top.cb_syn.char_path_n[89] ),
    .A1(\top.cb_syn.char_path_n[90] ),
    .A2(\top.cb_syn.char_path_n[93] ),
    .A3(\top.cb_syn.char_path_n[94] ),
    .S0(net498),
    .S1(net492),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04796_));
 sky130_fd_sc_hd__and2_1 _08577_ (.A(_02542_),
    .B(_04796_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04797_));
 sky130_fd_sc_hd__mux4_1 _08578_ (.A0(\top.cb_syn.char_path_n[91] ),
    .A1(\top.cb_syn.char_path_n[92] ),
    .A2(\top.cb_syn.char_path_n[95] ),
    .A3(\top.cb_syn.char_path_n[96] ),
    .S0(net498),
    .S1(net492),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04798_));
 sky130_fd_sc_hd__a21o_1 _08579_ (.A1(net496),
    .A2(_04798_),
    .B1(_02541_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04799_));
 sky130_fd_sc_hd__o221a_1 _08580_ (.A1(\top.cb_syn.end_cnt[3] ),
    .A2(_04795_),
    .B1(_04797_),
    .B2(_04799_),
    .C1(\top.cb_syn.end_cnt[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04800_));
 sky130_fd_sc_hd__mux4_1 _08581_ (.A0(\top.cb_syn.char_path_n[73] ),
    .A1(\top.cb_syn.char_path_n[74] ),
    .A2(\top.cb_syn.char_path_n[77] ),
    .A3(\top.cb_syn.char_path_n[78] ),
    .S0(net501),
    .S1(net495),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04801_));
 sky130_fd_sc_hd__and2_1 _08582_ (.A(_02542_),
    .B(_04801_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04802_));
 sky130_fd_sc_hd__mux4_1 _08583_ (.A0(\top.cb_syn.char_path_n[75] ),
    .A1(\top.cb_syn.char_path_n[76] ),
    .A2(\top.cb_syn.char_path_n[79] ),
    .A3(\top.cb_syn.char_path_n[80] ),
    .S0(net500),
    .S1(net494),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04803_));
 sky130_fd_sc_hd__a21o_1 _08584_ (.A1(net497),
    .A2(_04803_),
    .B1(_02541_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04804_));
 sky130_fd_sc_hd__mux4_1 _08585_ (.A0(\top.cb_syn.char_path_n[65] ),
    .A1(\top.cb_syn.char_path_n[66] ),
    .A2(\top.cb_syn.char_path_n[69] ),
    .A3(\top.cb_syn.char_path_n[70] ),
    .S0(net500),
    .S1(net494),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04805_));
 sky130_fd_sc_hd__mux4_1 _08586_ (.A0(\top.cb_syn.char_path_n[67] ),
    .A1(\top.cb_syn.char_path_n[68] ),
    .A2(\top.cb_syn.char_path_n[71] ),
    .A3(\top.cb_syn.char_path_n[72] ),
    .S0(net500),
    .S1(net494),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04806_));
 sky130_fd_sc_hd__mux2_1 _08587_ (.A0(_04805_),
    .A1(_04806_),
    .S(net497),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04807_));
 sky130_fd_sc_hd__o221a_1 _08588_ (.A1(_04802_),
    .A2(_04804_),
    .B1(_04807_),
    .B2(\top.cb_syn.end_cnt[3] ),
    .C1(_02540_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04808_));
 sky130_fd_sc_hd__or3_1 _08589_ (.A(\top.cb_syn.end_cnt[5] ),
    .B(_04800_),
    .C(_04808_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04809_));
 sky130_fd_sc_hd__mux4_1 _08590_ (.A0(\top.cb_syn.char_path_n[105] ),
    .A1(\top.cb_syn.char_path_n[106] ),
    .A2(\top.cb_syn.char_path_n[109] ),
    .A3(\top.cb_syn.char_path_n[110] ),
    .S0(net500),
    .S1(net494),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04810_));
 sky130_fd_sc_hd__and2_1 _08591_ (.A(_02542_),
    .B(_04810_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04811_));
 sky130_fd_sc_hd__mux4_1 _08592_ (.A0(\top.cb_syn.char_path_n[107] ),
    .A1(\top.cb_syn.char_path_n[108] ),
    .A2(\top.cb_syn.char_path_n[111] ),
    .A3(\top.cb_syn.char_path_n[112] ),
    .S0(net501),
    .S1(net495),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04812_));
 sky130_fd_sc_hd__a21o_1 _08593_ (.A1(net497),
    .A2(_04812_),
    .B1(_02541_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04813_));
 sky130_fd_sc_hd__mux4_1 _08594_ (.A0(\top.cb_syn.char_path_n[97] ),
    .A1(\top.cb_syn.char_path_n[98] ),
    .A2(\top.cb_syn.char_path_n[101] ),
    .A3(\top.cb_syn.char_path_n[102] ),
    .S0(net500),
    .S1(net494),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04814_));
 sky130_fd_sc_hd__mux4_1 _08595_ (.A0(\top.cb_syn.char_path_n[99] ),
    .A1(\top.cb_syn.char_path_n[100] ),
    .A2(\top.cb_syn.char_path_n[103] ),
    .A3(\top.cb_syn.char_path_n[104] ),
    .S0(net500),
    .S1(net494),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04815_));
 sky130_fd_sc_hd__mux2_1 _08596_ (.A0(_04814_),
    .A1(_04815_),
    .S(net497),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04816_));
 sky130_fd_sc_hd__o221a_1 _08597_ (.A1(_04811_),
    .A2(_04813_),
    .B1(_04816_),
    .B2(\top.cb_syn.end_cnt[3] ),
    .C1(_02540_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04817_));
 sky130_fd_sc_hd__mux4_1 _08598_ (.A0(\top.cb_syn.char_path_n[123] ),
    .A1(\top.cb_syn.char_path_n[124] ),
    .A2(\top.cb_syn.char_path_n[127] ),
    .A3(\top.cb_syn.curr_path[127] ),
    .S0(net498),
    .S1(net492),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04818_));
 sky130_fd_sc_hd__mux4_1 _08599_ (.A0(\top.cb_syn.char_path_n[121] ),
    .A1(\top.cb_syn.char_path_n[122] ),
    .A2(\top.cb_syn.char_path_n[125] ),
    .A3(\top.cb_syn.char_path_n[126] ),
    .S0(net498),
    .S1(net492),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04819_));
 sky130_fd_sc_hd__mux2_1 _08600_ (.A0(_04818_),
    .A1(_04819_),
    .S(_02542_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04820_));
 sky130_fd_sc_hd__mux4_1 _08601_ (.A0(\top.cb_syn.char_path_n[113] ),
    .A1(\top.cb_syn.char_path_n[114] ),
    .A2(\top.cb_syn.char_path_n[117] ),
    .A3(\top.cb_syn.char_path_n[118] ),
    .S0(net499),
    .S1(net493),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04821_));
 sky130_fd_sc_hd__and2_1 _08602_ (.A(_02542_),
    .B(_04821_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04822_));
 sky130_fd_sc_hd__mux4_1 _08603_ (.A0(\top.cb_syn.char_path_n[115] ),
    .A1(\top.cb_syn.char_path_n[116] ),
    .A2(\top.cb_syn.char_path_n[119] ),
    .A3(\top.cb_syn.char_path_n[120] ),
    .S0(net499),
    .S1(net493),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04823_));
 sky130_fd_sc_hd__a21o_1 _08604_ (.A1(net496),
    .A2(_04823_),
    .B1(\top.cb_syn.end_cnt[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04824_));
 sky130_fd_sc_hd__o221a_1 _08605_ (.A1(_02541_),
    .A2(_04820_),
    .B1(_04822_),
    .B2(_04824_),
    .C1(\top.cb_syn.end_cnt[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04825_));
 sky130_fd_sc_hd__or3b_1 _08606_ (.A(_04817_),
    .B(_04825_),
    .C_N(\top.cb_syn.end_cnt[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04826_));
 sky130_fd_sc_hd__mux4_1 _08607_ (.A0(\top.cb_syn.char_path_n[25] ),
    .A1(\top.cb_syn.char_path_n[26] ),
    .A2(\top.cb_syn.char_path_n[29] ),
    .A3(\top.cb_syn.char_path_n[30] ),
    .S0(net498),
    .S1(net492),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04827_));
 sky130_fd_sc_hd__mux4_1 _08608_ (.A0(\top.cb_syn.char_path_n[27] ),
    .A1(\top.cb_syn.char_path_n[28] ),
    .A2(\top.cb_syn.char_path_n[31] ),
    .A3(\top.cb_syn.char_path_n[32] ),
    .S0(net498),
    .S1(net492),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04828_));
 sky130_fd_sc_hd__a21o_1 _08609_ (.A1(net496),
    .A2(_04828_),
    .B1(_02541_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04829_));
 sky130_fd_sc_hd__a21o_1 _08610_ (.A1(_02542_),
    .A2(_04827_),
    .B1(_04829_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04830_));
 sky130_fd_sc_hd__mux4_1 _08611_ (.A0(\top.cb_syn.char_path_n[17] ),
    .A1(\top.cb_syn.char_path_n[18] ),
    .A2(\top.cb_syn.char_path_n[21] ),
    .A3(\top.cb_syn.char_path_n[22] ),
    .S0(net499),
    .S1(net493),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04831_));
 sky130_fd_sc_hd__mux4_1 _08612_ (.A0(\top.cb_syn.char_path_n[19] ),
    .A1(\top.cb_syn.char_path_n[20] ),
    .A2(\top.cb_syn.char_path_n[23] ),
    .A3(\top.cb_syn.char_path_n[24] ),
    .S0(net499),
    .S1(net493),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04832_));
 sky130_fd_sc_hd__mux2_1 _08613_ (.A0(_04831_),
    .A1(_04832_),
    .S(net496),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04833_));
 sky130_fd_sc_hd__o211a_1 _08614_ (.A1(\top.cb_syn.end_cnt[3] ),
    .A2(_04833_),
    .B1(_04830_),
    .C1(\top.cb_syn.end_cnt[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04834_));
 sky130_fd_sc_hd__mux4_1 _08615_ (.A0(\top.cb_syn.char_path_n[11] ),
    .A1(\top.cb_syn.char_path_n[12] ),
    .A2(\top.cb_syn.char_path_n[15] ),
    .A3(\top.cb_syn.char_path_n[16] ),
    .S0(net501),
    .S1(net495),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04835_));
 sky130_fd_sc_hd__mux4_1 _08616_ (.A0(\top.cb_syn.char_path_n[9] ),
    .A1(\top.cb_syn.char_path_n[10] ),
    .A2(\top.cb_syn.char_path_n[13] ),
    .A3(\top.cb_syn.char_path_n[14] ),
    .S0(net501),
    .S1(net495),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04836_));
 sky130_fd_sc_hd__mux2_1 _08617_ (.A0(_04835_),
    .A1(_04836_),
    .S(_02542_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04837_));
 sky130_fd_sc_hd__or2_1 _08618_ (.A(_02541_),
    .B(_04837_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04838_));
 sky130_fd_sc_hd__mux4_1 _08619_ (.A0(\top.cb_syn.char_path_n[1] ),
    .A1(\top.cb_syn.char_path_n[2] ),
    .A2(\top.cb_syn.char_path_n[5] ),
    .A3(\top.cb_syn.char_path_n[6] ),
    .S0(net501),
    .S1(net495),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04839_));
 sky130_fd_sc_hd__mux4_1 _08620_ (.A0(\top.cb_syn.char_path_n[3] ),
    .A1(\top.cb_syn.char_path_n[4] ),
    .A2(\top.cb_syn.char_path_n[7] ),
    .A3(\top.cb_syn.char_path_n[8] ),
    .S0(net501),
    .S1(net495),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04840_));
 sky130_fd_sc_hd__mux2_1 _08621_ (.A0(_04839_),
    .A1(_04840_),
    .S(net497),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04841_));
 sky130_fd_sc_hd__or2_1 _08622_ (.A(\top.cb_syn.end_cnt[3] ),
    .B(_04841_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04842_));
 sky130_fd_sc_hd__a311o_1 _08623_ (.A1(_02540_),
    .A2(_04838_),
    .A3(_04842_),
    .B1(_04834_),
    .C1(\top.cb_syn.end_cnt[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04843_));
 sky130_fd_sc_hd__mux4_1 _08624_ (.A0(\top.cb_syn.char_path_n[59] ),
    .A1(\top.cb_syn.char_path_n[60] ),
    .A2(\top.cb_syn.char_path_n[63] ),
    .A3(\top.cb_syn.char_path_n[64] ),
    .S0(net498),
    .S1(net492),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04844_));
 sky130_fd_sc_hd__mux4_1 _08625_ (.A0(\top.cb_syn.char_path_n[57] ),
    .A1(\top.cb_syn.char_path_n[58] ),
    .A2(\top.cb_syn.char_path_n[61] ),
    .A3(\top.cb_syn.char_path_n[62] ),
    .S0(net498),
    .S1(net492),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04845_));
 sky130_fd_sc_hd__mux2_1 _08626_ (.A0(_04844_),
    .A1(_04845_),
    .S(_02542_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04846_));
 sky130_fd_sc_hd__mux4_1 _08627_ (.A0(\top.cb_syn.char_path_n[49] ),
    .A1(\top.cb_syn.char_path_n[50] ),
    .A2(\top.cb_syn.char_path_n[53] ),
    .A3(\top.cb_syn.char_path_n[54] ),
    .S0(net499),
    .S1(net493),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04847_));
 sky130_fd_sc_hd__mux4_1 _08628_ (.A0(\top.cb_syn.char_path_n[51] ),
    .A1(\top.cb_syn.char_path_n[52] ),
    .A2(\top.cb_syn.char_path_n[55] ),
    .A3(\top.cb_syn.char_path_n[56] ),
    .S0(net499),
    .S1(net493),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04848_));
 sky130_fd_sc_hd__mux2_1 _08629_ (.A0(_04847_),
    .A1(_04848_),
    .S(net496),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04849_));
 sky130_fd_sc_hd__mux2_1 _08630_ (.A0(_04846_),
    .A1(_04849_),
    .S(_02541_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04850_));
 sky130_fd_sc_hd__mux4_1 _08631_ (.A0(\top.cb_syn.char_path_n[41] ),
    .A1(\top.cb_syn.char_path_n[42] ),
    .A2(\top.cb_syn.char_path_n[45] ),
    .A3(\top.cb_syn.char_path_n[46] ),
    .S0(net500),
    .S1(net494),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04851_));
 sky130_fd_sc_hd__mux4_1 _08632_ (.A0(\top.cb_syn.char_path_n[43] ),
    .A1(\top.cb_syn.char_path_n[44] ),
    .A2(\top.cb_syn.char_path_n[47] ),
    .A3(\top.cb_syn.char_path_n[48] ),
    .S0(net500),
    .S1(net494),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04852_));
 sky130_fd_sc_hd__and2_1 _08633_ (.A(net497),
    .B(_04852_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04853_));
 sky130_fd_sc_hd__a211o_1 _08634_ (.A1(_02542_),
    .A2(_04851_),
    .B1(_04853_),
    .C1(_02541_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04854_));
 sky130_fd_sc_hd__mux4_1 _08635_ (.A0(\top.cb_syn.char_path_n[33] ),
    .A1(\top.cb_syn.char_path_n[34] ),
    .A2(\top.cb_syn.char_path_n[37] ),
    .A3(\top.cb_syn.char_path_n[38] ),
    .S0(net500),
    .S1(net494),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04855_));
 sky130_fd_sc_hd__mux4_1 _08636_ (.A0(\top.cb_syn.char_path_n[35] ),
    .A1(\top.cb_syn.char_path_n[36] ),
    .A2(\top.cb_syn.char_path_n[39] ),
    .A3(\top.cb_syn.char_path_n[40] ),
    .S0(net500),
    .S1(net494),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04856_));
 sky130_fd_sc_hd__mux2_1 _08637_ (.A0(_04855_),
    .A1(_04856_),
    .S(net497),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04857_));
 sky130_fd_sc_hd__o211a_1 _08638_ (.A1(\top.cb_syn.end_cnt[3] ),
    .A2(_04857_),
    .B1(_04854_),
    .C1(_02540_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04858_));
 sky130_fd_sc_hd__a21oi_1 _08639_ (.A1(\top.cb_syn.end_cnt[4] ),
    .A2(_04850_),
    .B1(_04858_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04859_));
 sky130_fd_sc_hd__a21oi_1 _08640_ (.A1(\top.cb_syn.end_cnt[5] ),
    .A2(_04859_),
    .B1(\top.cb_syn.end_cnt[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04860_));
 sky130_fd_sc_hd__a32o_1 _08641_ (.A1(\top.cb_syn.end_cnt[6] ),
    .A2(_04809_),
    .A3(_04826_),
    .B1(_04843_),
    .B2(_04860_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04861_));
 sky130_fd_sc_hd__and2b_1 _08642_ (.A_N(_04792_),
    .B(_04861_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04862_));
 sky130_fd_sc_hd__o21ai_1 _08643_ (.A1(net520),
    .A2(\top.cb_syn.curr_state[5] ),
    .B1(_04770_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04863_));
 sky130_fd_sc_hd__or3b_1 _08644_ (.A(_04862_),
    .B(_04863_),
    .C_N(\top.cb_syn.cb_enable ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04864_));
 sky130_fd_sc_hd__a22o_1 _08645_ (.A1(net519),
    .A2(_04770_),
    .B1(_04864_),
    .B2(net1647),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01480_));
 sky130_fd_sc_hd__or3_1 _08646_ (.A(_04196_),
    .B(_04768_),
    .C(_04769_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04865_));
 sky130_fd_sc_hd__mux2_1 _08647_ (.A0(net519),
    .A1(net1037),
    .S(_04865_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01479_));
 sky130_fd_sc_hd__or2_2 _08648_ (.A(_02888_),
    .B(_04863_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04866_));
 sky130_fd_sc_hd__a21oi_1 _08649_ (.A1(_02538_),
    .A2(_04791_),
    .B1(_04866_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04867_));
 sky130_fd_sc_hd__or2_2 _08650_ (.A(net520),
    .B(_04866_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04868_));
 sky130_fd_sc_hd__or2_1 _08651_ (.A(_04791_),
    .B(_04868_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04869_));
 sky130_fd_sc_hd__mux2_1 _08652_ (.A0(_04867_),
    .A1(_04869_),
    .S(\top.cb_syn.end_cnt[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01478_));
 sky130_fd_sc_hd__o31a_1 _08653_ (.A1(\top.cb_syn.end_cnt[4] ),
    .A2(_04790_),
    .A3(_04866_),
    .B1(\top.cb_syn.end_cnt[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04870_));
 sky130_fd_sc_hd__or2_1 _08654_ (.A(_04867_),
    .B(_04870_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01477_));
 sky130_fd_sc_hd__a21oi_1 _08655_ (.A1(_02538_),
    .A2(_04790_),
    .B1(_04866_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04871_));
 sky130_fd_sc_hd__or2_1 _08656_ (.A(_02540_),
    .B(_04790_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04872_));
 sky130_fd_sc_hd__o22a_1 _08657_ (.A1(\top.cb_syn.end_cnt[4] ),
    .A2(_04871_),
    .B1(_04872_),
    .B2(_04868_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01476_));
 sky130_fd_sc_hd__or3b_1 _08658_ (.A(_04866_),
    .B(net493),
    .C_N(_04789_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04873_));
 sky130_fd_sc_hd__a21o_1 _08659_ (.A1(\top.cb_syn.end_cnt[3] ),
    .A2(_04873_),
    .B1(_04871_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01475_));
 sky130_fd_sc_hd__o21ba_1 _08660_ (.A1(\top.cb_syn.char_path_n[0] ),
    .A2(_04789_),
    .B1_N(_04866_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04874_));
 sky130_fd_sc_hd__nand2_1 _08661_ (.A(net492),
    .B(_04789_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04875_));
 sky130_fd_sc_hd__o22a_1 _08662_ (.A1(net492),
    .A2(_04874_),
    .B1(_04875_),
    .B2(_04868_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01474_));
 sky130_fd_sc_hd__or2_1 _08663_ (.A(net499),
    .B(_04866_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04876_));
 sky130_fd_sc_hd__a21o_1 _08664_ (.A1(net496),
    .A2(_04876_),
    .B1(_04874_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01473_));
 sky130_fd_sc_hd__a21bo_1 _08665_ (.A1(net499),
    .A2(_04868_),
    .B1_N(_04876_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01472_));
 sky130_fd_sc_hd__a21oi_1 _08666_ (.A1(\top.cb_syn.cb_enable ),
    .A2(_04792_),
    .B1(_04868_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04877_));
 sky130_fd_sc_hd__a22o_1 _08667_ (.A1(net1621),
    .A2(_04866_),
    .B1(_04877_),
    .B2(_04861_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01471_));
 sky130_fd_sc_hd__o221ai_2 _08668_ (.A1(net522),
    .A2(net523),
    .B1(_04189_),
    .B2(_04190_),
    .C1(_04561_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04878_));
 sky130_fd_sc_hd__or2_2 _08669_ (.A(_04605_),
    .B(_04878_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04879_));
 sky130_fd_sc_hd__nand2_1 _08670_ (.A(\top.cb_syn.i[1] ),
    .B(\top.cb_syn.i[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04880_));
 sky130_fd_sc_hd__and4_1 _08671_ (.A(\top.cb_syn.i[3] ),
    .B(\top.cb_syn.i[2] ),
    .C(\top.cb_syn.i[1] ),
    .D(\top.cb_syn.i[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04881_));
 sky130_fd_sc_hd__inv_2 _08672_ (.A(_04881_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04882_));
 sky130_fd_sc_hd__nand2_1 _08673_ (.A(\top.cb_syn.i[4] ),
    .B(_04881_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04883_));
 sky130_fd_sc_hd__and3_1 _08674_ (.A(\top.cb_syn.i[5] ),
    .B(\top.cb_syn.i[4] ),
    .C(_04881_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04884_));
 sky130_fd_sc_hd__o21bai_1 _08675_ (.A1(\top.cb_syn.curr_state[2] ),
    .A2(_04884_),
    .B1_N(_04879_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04885_));
 sky130_fd_sc_hd__nor2_1 _08676_ (.A(\top.cb_syn.curr_state[2] ),
    .B(_04878_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04886_));
 sky130_fd_sc_hd__and2_1 _08677_ (.A(_04884_),
    .B(_04886_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04887_));
 sky130_fd_sc_hd__mux2_1 _08678_ (.A0(_04887_),
    .A1(_04885_),
    .S(net1649),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01470_));
 sky130_fd_sc_hd__nor2_1 _08679_ (.A(_04879_),
    .B(_04883_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04888_));
 sky130_fd_sc_hd__o21a_1 _08680_ (.A1(net1622),
    .A2(_04888_),
    .B1(_04885_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01469_));
 sky130_fd_sc_hd__or2_1 _08681_ (.A(\top.cb_syn.i[4] ),
    .B(_04881_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04889_));
 sky130_fd_sc_hd__a32o_1 _08682_ (.A1(_04883_),
    .A2(_04886_),
    .A3(_04889_),
    .B1(_04879_),
    .B2(net1783),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01468_));
 sky130_fd_sc_hd__a31o_1 _08683_ (.A1(\top.cb_syn.i[2] ),
    .A2(\top.cb_syn.i[1] ),
    .A3(\top.cb_syn.i[0] ),
    .B1(\top.cb_syn.i[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04890_));
 sky130_fd_sc_hd__a32o_1 _08684_ (.A1(_04882_),
    .A2(_04886_),
    .A3(_04890_),
    .B1(_04879_),
    .B2(net1714),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01467_));
 sky130_fd_sc_hd__xnor2_1 _08685_ (.A(\top.cb_syn.i[2] ),
    .B(_04880_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04891_));
 sky130_fd_sc_hd__a22o_1 _08686_ (.A1(\top.cb_syn.i[2] ),
    .A2(_04879_),
    .B1(_04886_),
    .B2(_04891_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01466_));
 sky130_fd_sc_hd__or2_1 _08687_ (.A(\top.cb_syn.i[1] ),
    .B(\top.cb_syn.i[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04892_));
 sky130_fd_sc_hd__a32o_1 _08688_ (.A1(_04880_),
    .A2(_04886_),
    .A3(_04892_),
    .B1(_04879_),
    .B2(net1688),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01465_));
 sky130_fd_sc_hd__mux2_1 _08689_ (.A0(_04886_),
    .A1(_04879_),
    .S(\top.cb_syn.i[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01464_));
 sky130_fd_sc_hd__and4_1 _08690_ (.A(\top.cb_syn.cb_enable ),
    .B(\top.cb_syn.curr_state[5] ),
    .C(net464),
    .D(_04792_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04893_));
 sky130_fd_sc_hd__a31o_1 _08691_ (.A1(\top.cb_syn.end_check ),
    .A2(_04861_),
    .A3(_04893_),
    .B1(net1482),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01463_));
 sky130_fd_sc_hd__o211ai_1 _08692_ (.A1(_02543_),
    .A2(_04562_),
    .B1(_04208_),
    .C1(_04179_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04894_));
 sky130_fd_sc_hd__a32o_1 _08693_ (.A1(net515),
    .A2(_04208_),
    .A3(_04562_),
    .B1(_04894_),
    .B2(net1572),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01462_));
 sky130_fd_sc_hd__a21oi_1 _08694_ (.A1(_02566_),
    .A2(\top.header_synthesis.start ),
    .B1(_03389_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04895_));
 sky130_fd_sc_hd__nor2_1 _08695_ (.A(_02544_),
    .B(_03389_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04896_));
 sky130_fd_sc_hd__and4_1 _08696_ (.A(\top.header_synthesis.count[4] ),
    .B(\top.header_synthesis.count[3] ),
    .C(\top.header_synthesis.count[2] ),
    .D(\top.header_synthesis.count[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04897_));
 sky130_fd_sc_hd__and2_1 _08697_ (.A(\top.header_synthesis.count[1] ),
    .B(_04896_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04898_));
 sky130_fd_sc_hd__and3_1 _08698_ (.A(\top.header_synthesis.count[2] ),
    .B(\top.header_synthesis.count[1] ),
    .C(_04896_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04899_));
 sky130_fd_sc_hd__and3_1 _08699_ (.A(\top.header_synthesis.count[3] ),
    .B(\top.header_synthesis.count[2] ),
    .C(_04898_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04900_));
 sky130_fd_sc_hd__a21oi_1 _08700_ (.A1(_04896_),
    .A2(_04897_),
    .B1(_04895_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04901_));
 sky130_fd_sc_hd__and3_1 _08701_ (.A(\top.header_synthesis.count[5] ),
    .B(_04896_),
    .C(_04897_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04902_));
 sky130_fd_sc_hd__a21oi_1 _08702_ (.A1(\top.header_synthesis.count[6] ),
    .A2(_04902_),
    .B1(_04895_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04903_));
 sky130_fd_sc_hd__and4_1 _08703_ (.A(\top.header_synthesis.count[0] ),
    .B(_02566_),
    .C(_03370_),
    .D(_04897_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04904_));
 sky130_fd_sc_hd__and4b_1 _08704_ (.A_N(\top.header_synthesis.count[7] ),
    .B(\top.header_synthesis.count[6] ),
    .C(\top.header_synthesis.count[5] ),
    .D(_04904_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04905_));
 sky130_fd_sc_hd__a21o_1 _08705_ (.A1(net1430),
    .A2(_04903_),
    .B1(_04905_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01461_));
 sky130_fd_sc_hd__o21a_1 _08706_ (.A1(net1652),
    .A2(_04902_),
    .B1(_04903_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01460_));
 sky130_fd_sc_hd__mux2_1 _08707_ (.A0(_04904_),
    .A1(_04901_),
    .S(net1739),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01459_));
 sky130_fd_sc_hd__o21a_1 _08708_ (.A1(net1508),
    .A2(_04900_),
    .B1(_04901_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01458_));
 sky130_fd_sc_hd__a21o_1 _08709_ (.A1(\top.header_synthesis.enable ),
    .A2(\top.header_synthesis.char_added ),
    .B1(\top.header_synthesis.write_num_lefts ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04906_));
 sky130_fd_sc_hd__a21bo_1 _08710_ (.A1(_03375_),
    .A2(_04906_),
    .B1_N(_04895_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04907_));
 sky130_fd_sc_hd__o21ai_1 _08711_ (.A1(\top.header_synthesis.count[3] ),
    .A2(_04899_),
    .B1(_04907_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04908_));
 sky130_fd_sc_hd__nor2_1 _08712_ (.A(_04900_),
    .B(_04908_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_01457_));
 sky130_fd_sc_hd__o21ai_1 _08713_ (.A1(\top.header_synthesis.count[2] ),
    .A2(_04898_),
    .B1(_04907_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04909_));
 sky130_fd_sc_hd__nor2_1 _08714_ (.A(_04899_),
    .B(_04909_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_01456_));
 sky130_fd_sc_hd__o21ai_1 _08715_ (.A1(\top.header_synthesis.count[1] ),
    .A2(_04896_),
    .B1(_04907_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04910_));
 sky130_fd_sc_hd__nor2_1 _08716_ (.A(_04898_),
    .B(_04910_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_01455_));
 sky130_fd_sc_hd__nand2_1 _08717_ (.A(_02544_),
    .B(_03389_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04911_));
 sky130_fd_sc_hd__and3b_1 _08718_ (.A_N(_04896_),
    .B(_04907_),
    .C(_04911_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01454_));
 sky130_fd_sc_hd__o21a_1 _08719_ (.A1(net431),
    .A2(_04255_),
    .B1(net980),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01453_));
 sky130_fd_sc_hd__nor2_1 _08720_ (.A(net542),
    .B(_02591_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04912_));
 sky130_fd_sc_hd__nor2_1 _08721_ (.A(net304),
    .B(_04912_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04913_));
 sky130_fd_sc_hd__a21boi_1 _08722_ (.A1(\top.sram_interface.TRN_counter[1] ),
    .A2(\top.sram_interface.TRN_counter[0] ),
    .B1_N(\top.sram_interface.TRN_counter[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04914_));
 sky130_fd_sc_hd__o21a_1 _08723_ (.A1(_02913_),
    .A2(_04914_),
    .B1(_02589_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04915_));
 sky130_fd_sc_hd__mux2_1 _08724_ (.A0(_04915_),
    .A1(\top.sram_interface.TRN_counter[2] ),
    .S(_04913_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01452_));
 sky130_fd_sc_hd__nand2b_1 _08725_ (.A_N(_04913_),
    .B(\top.sram_interface.TRN_counter[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04916_));
 sky130_fd_sc_hd__xnor2_1 _08726_ (.A(net1678),
    .B(_04916_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_01451_));
 sky130_fd_sc_hd__o21a_1 _08727_ (.A1(\top.sram_interface.TRN_counter[0] ),
    .A2(_04912_),
    .B1(_04916_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01450_));
 sky130_fd_sc_hd__nand2_2 _08728_ (.A(net425),
    .B(net508),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04917_));
 sky130_fd_sc_hd__mux4_1 _08729_ (.A0(\top.path[56] ),
    .A1(\top.path[57] ),
    .A2(\top.path[58] ),
    .A3(\top.path[59] ),
    .S0(net508),
    .S1(net506),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04918_));
 sky130_fd_sc_hd__mux2_1 _08730_ (.A0(\top.path[62] ),
    .A1(\top.path[63] ),
    .S(net511),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04919_));
 sky130_fd_sc_hd__or2_1 _08731_ (.A(net426),
    .B(_04919_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04920_));
 sky130_fd_sc_hd__o221a_1 _08732_ (.A1(\top.path[60] ),
    .A2(net404),
    .B1(net324),
    .B2(\top.path[61] ),
    .C1(net505),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04921_));
 sky130_fd_sc_hd__a22o_1 _08733_ (.A1(net430),
    .A2(_04918_),
    .B1(_04920_),
    .B2(_04921_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04922_));
 sky130_fd_sc_hd__mux2_1 _08734_ (.A0(\top.path[50] ),
    .A1(\top.path[51] ),
    .S(net511),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04923_));
 sky130_fd_sc_hd__or2_1 _08735_ (.A(net426),
    .B(_04923_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04924_));
 sky130_fd_sc_hd__o221a_1 _08736_ (.A1(\top.path[48] ),
    .A2(net404),
    .B1(net324),
    .B2(\top.path[49] ),
    .C1(net429),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04925_));
 sky130_fd_sc_hd__mux4_1 _08737_ (.A0(\top.path[52] ),
    .A1(\top.path[53] ),
    .A2(\top.path[54] ),
    .A3(\top.path[55] ),
    .S0(net511),
    .S1(net507),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04926_));
 sky130_fd_sc_hd__mux2_1 _08738_ (.A0(\top.path[126] ),
    .A1(\top.path[127] ),
    .S(net511),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04927_));
 sky130_fd_sc_hd__o221a_1 _08739_ (.A1(\top.path[125] ),
    .A2(net324),
    .B1(_04927_),
    .B2(net427),
    .C1(net505),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04928_));
 sky130_fd_sc_hd__o21a_1 _08740_ (.A1(\top.path[124] ),
    .A2(net405),
    .B1(_04928_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04929_));
 sky130_fd_sc_hd__mux2_1 _08741_ (.A0(\top.path[122] ),
    .A1(\top.path[123] ),
    .S(net512),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04930_));
 sky130_fd_sc_hd__o221a_1 _08742_ (.A1(\top.path[120] ),
    .A2(net403),
    .B1(net323),
    .B2(\top.path[121] ),
    .C1(net429),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04931_));
 sky130_fd_sc_hd__o21a_1 _08743_ (.A1(net425),
    .A2(_04930_),
    .B1(_04931_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04932_));
 sky130_fd_sc_hd__mux2_1 _08744_ (.A0(\top.path[118] ),
    .A1(\top.path[119] ),
    .S(net512),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04933_));
 sky130_fd_sc_hd__or2_1 _08745_ (.A(net428),
    .B(_04933_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04934_));
 sky130_fd_sc_hd__o221a_1 _08746_ (.A1(\top.path[116] ),
    .A2(net403),
    .B1(net323),
    .B2(\top.path[117] ),
    .C1(net505),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04935_));
 sky130_fd_sc_hd__mux4_1 _08747_ (.A0(\top.path[112] ),
    .A1(\top.path[113] ),
    .A2(\top.path[114] ),
    .A3(\top.path[115] ),
    .S0(net508),
    .S1(net506),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04936_));
 sky130_fd_sc_hd__mux2_1 _08748_ (.A0(\top.path[26] ),
    .A1(\top.path[27] ),
    .S(net509),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04937_));
 sky130_fd_sc_hd__or2_1 _08749_ (.A(net425),
    .B(_04937_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04938_));
 sky130_fd_sc_hd__mux2_1 _08750_ (.A0(\top.path[18] ),
    .A1(\top.path[19] ),
    .S(net508),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04939_));
 sky130_fd_sc_hd__or2_1 _08751_ (.A(net425),
    .B(_04939_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04940_));
 sky130_fd_sc_hd__mux2_1 _08752_ (.A0(\top.path[30] ),
    .A1(\top.path[31] ),
    .S(net511),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04941_));
 sky130_fd_sc_hd__o221a_1 _08753_ (.A1(\top.path[29] ),
    .A2(net325),
    .B1(_04941_),
    .B2(net427),
    .C1(net502),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04942_));
 sky130_fd_sc_hd__o21a_1 _08754_ (.A1(\top.path[28] ),
    .A2(net405),
    .B1(_04942_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04943_));
 sky130_fd_sc_hd__mux2_1 _08755_ (.A0(\top.path[22] ),
    .A1(\top.path[23] ),
    .S(net512),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04944_));
 sky130_fd_sc_hd__o221a_1 _08756_ (.A1(\top.path[20] ),
    .A2(net403),
    .B1(net323),
    .B2(\top.path[21] ),
    .C1(_02547_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04945_));
 sky130_fd_sc_hd__o21a_1 _08757_ (.A1(net428),
    .A2(_04944_),
    .B1(_04945_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04946_));
 sky130_fd_sc_hd__mux2_1 _08758_ (.A0(\top.path[86] ),
    .A1(\top.path[87] ),
    .S(net508),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04947_));
 sky130_fd_sc_hd__or2_1 _08759_ (.A(net425),
    .B(_04947_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04948_));
 sky130_fd_sc_hd__o221a_1 _08760_ (.A1(\top.path[84] ),
    .A2(net402),
    .B1(net323),
    .B2(\top.path[85] ),
    .C1(net504),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04949_));
 sky130_fd_sc_hd__mux4_1 _08761_ (.A0(\top.path[80] ),
    .A1(\top.path[81] ),
    .A2(\top.path[82] ),
    .A3(\top.path[83] ),
    .S0(net508),
    .S1(net506),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04950_));
 sky130_fd_sc_hd__mux2_1 _08762_ (.A0(\top.path[94] ),
    .A1(\top.path[95] ),
    .S(net511),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04951_));
 sky130_fd_sc_hd__o221a_1 _08763_ (.A1(\top.path[93] ),
    .A2(net323),
    .B1(_04951_),
    .B2(net425),
    .C1(net504),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04952_));
 sky130_fd_sc_hd__o21a_1 _08764_ (.A1(\top.path[92] ),
    .A2(net402),
    .B1(_04952_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04953_));
 sky130_fd_sc_hd__mux2_1 _08765_ (.A0(\top.path[90] ),
    .A1(\top.path[91] ),
    .S(net508),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04954_));
 sky130_fd_sc_hd__o221a_1 _08766_ (.A1(\top.path[88] ),
    .A2(net402),
    .B1(net323),
    .B2(\top.path[89] ),
    .C1(net429),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04955_));
 sky130_fd_sc_hd__o21a_1 _08767_ (.A1(net425),
    .A2(_04954_),
    .B1(_04955_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04956_));
 sky130_fd_sc_hd__or3_1 _08768_ (.A(_02547_),
    .B(_04929_),
    .C(_04932_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04957_));
 sky130_fd_sc_hd__a221o_1 _08769_ (.A1(_04934_),
    .A2(_04935_),
    .B1(_04936_),
    .B2(net429),
    .C1(net502),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04958_));
 sky130_fd_sc_hd__or3_1 _08770_ (.A(_02547_),
    .B(_04953_),
    .C(_04956_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04959_));
 sky130_fd_sc_hd__a221o_1 _08771_ (.A1(_04948_),
    .A2(_04949_),
    .B1(_04950_),
    .B2(net429),
    .C1(net502),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04960_));
 sky130_fd_sc_hd__a31o_1 _08772_ (.A1(_02546_),
    .A2(_04959_),
    .A3(_04960_),
    .B1(_02545_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04961_));
 sky130_fd_sc_hd__a31o_1 _08773_ (.A1(\top.translation.index[5] ),
    .A2(_04957_),
    .A3(_04958_),
    .B1(_04961_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04962_));
 sky130_fd_sc_hd__or3_1 _08774_ (.A(net430),
    .B(_04943_),
    .C(_04946_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04963_));
 sky130_fd_sc_hd__o221a_1 _08775_ (.A1(\top.path[24] ),
    .A2(net402),
    .B1(net323),
    .B2(\top.path[25] ),
    .C1(net502),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04964_));
 sky130_fd_sc_hd__o221a_1 _08776_ (.A1(\top.path[16] ),
    .A2(net403),
    .B1(_04917_),
    .B2(\top.path[17] ),
    .C1(_02547_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04965_));
 sky130_fd_sc_hd__a221o_1 _08777_ (.A1(_04938_),
    .A2(_04964_),
    .B1(_04965_),
    .B2(_04940_),
    .C1(net504),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04966_));
 sky130_fd_sc_hd__a221o_1 _08778_ (.A1(_04924_),
    .A2(_04925_),
    .B1(_04926_),
    .B2(net505),
    .C1(net503),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04967_));
 sky130_fd_sc_hd__o211a_1 _08779_ (.A1(_02547_),
    .A2(_04922_),
    .B1(_04967_),
    .C1(\top.translation.index[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04968_));
 sky130_fd_sc_hd__a311o_1 _08780_ (.A1(_02546_),
    .A2(_04963_),
    .A3(_04966_),
    .B1(_04968_),
    .C1(\top.translation.index[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04969_));
 sky130_fd_sc_hd__mux2_1 _08781_ (.A0(\top.path[14] ),
    .A1(\top.path[15] ),
    .S(net510),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04970_));
 sky130_fd_sc_hd__or2_1 _08782_ (.A(net426),
    .B(_04970_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04971_));
 sky130_fd_sc_hd__o221a_1 _08783_ (.A1(\top.path[12] ),
    .A2(net404),
    .B1(net324),
    .B2(\top.path[13] ),
    .C1(\top.translation.index[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04972_));
 sky130_fd_sc_hd__mux2_1 _08784_ (.A0(\top.path[10] ),
    .A1(\top.path[11] ),
    .S(net510),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04973_));
 sky130_fd_sc_hd__or2_1 _08785_ (.A(\top.path[8] ),
    .B(net404),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04974_));
 sky130_fd_sc_hd__o221a_1 _08786_ (.A1(\top.path[9] ),
    .A2(net324),
    .B1(_04973_),
    .B2(net426),
    .C1(net429),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04975_));
 sky130_fd_sc_hd__a22o_1 _08787_ (.A1(_04971_),
    .A2(_04972_),
    .B1(_04974_),
    .B2(_04975_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04976_));
 sky130_fd_sc_hd__mux4_1 _08788_ (.A0(\top.path[4] ),
    .A1(\top.path[5] ),
    .A2(\top.path[6] ),
    .A3(\top.path[7] ),
    .S0(net510),
    .S1(net507),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04977_));
 sky130_fd_sc_hd__mux2_1 _08789_ (.A0(\top.path[2] ),
    .A1(\top.path[3] ),
    .S(net510),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04978_));
 sky130_fd_sc_hd__o221a_1 _08790_ (.A1(\top.path[0] ),
    .A2(net404),
    .B1(net324),
    .B2(\top.path[1] ),
    .C1(net429),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04979_));
 sky130_fd_sc_hd__o21a_1 _08791_ (.A1(net426),
    .A2(_04978_),
    .B1(_04979_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04980_));
 sky130_fd_sc_hd__a21o_1 _08792_ (.A1(\top.translation.index[2] ),
    .A2(_04977_),
    .B1(net503),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04981_));
 sky130_fd_sc_hd__o22a_1 _08793_ (.A1(_02547_),
    .A2(_04976_),
    .B1(_04980_),
    .B2(_04981_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04982_));
 sky130_fd_sc_hd__mux2_1 _08794_ (.A0(\top.path[78] ),
    .A1(\top.path[79] ),
    .S(net511),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04983_));
 sky130_fd_sc_hd__o221a_1 _08795_ (.A1(\top.path[76] ),
    .A2(net404),
    .B1(net324),
    .B2(\top.path[77] ),
    .C1(net503),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04984_));
 sky130_fd_sc_hd__o21a_1 _08796_ (.A1(net426),
    .A2(_04983_),
    .B1(_04984_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04985_));
 sky130_fd_sc_hd__mux2_1 _08797_ (.A0(\top.path[70] ),
    .A1(\top.path[71] ),
    .S(net510),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04986_));
 sky130_fd_sc_hd__o221a_1 _08798_ (.A1(\top.path[69] ),
    .A2(net324),
    .B1(_04986_),
    .B2(net426),
    .C1(_02547_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04987_));
 sky130_fd_sc_hd__o21a_1 _08799_ (.A1(\top.path[68] ),
    .A2(net404),
    .B1(_04987_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04988_));
 sky130_fd_sc_hd__mux2_1 _08800_ (.A0(\top.path[66] ),
    .A1(\top.path[67] ),
    .S(net510),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04989_));
 sky130_fd_sc_hd__or2_1 _08801_ (.A(net426),
    .B(_04989_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04990_));
 sky130_fd_sc_hd__o221a_1 _08802_ (.A1(\top.path[64] ),
    .A2(net404),
    .B1(net324),
    .B2(\top.path[65] ),
    .C1(_02547_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04991_));
 sky130_fd_sc_hd__mux4_1 _08803_ (.A0(\top.path[72] ),
    .A1(\top.path[73] ),
    .A2(\top.path[74] ),
    .A3(\top.path[75] ),
    .S0(net511),
    .S1(net507),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04992_));
 sky130_fd_sc_hd__a221o_1 _08804_ (.A1(_04990_),
    .A2(_04991_),
    .B1(_04992_),
    .B2(net503),
    .C1(\top.translation.index[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04993_));
 sky130_fd_sc_hd__mux2_1 _08805_ (.A0(\top.path[46] ),
    .A1(\top.path[47] ),
    .S(net510),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04994_));
 sky130_fd_sc_hd__o221a_1 _08806_ (.A1(\top.path[44] ),
    .A2(net404),
    .B1(net324),
    .B2(\top.path[45] ),
    .C1(net505),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04995_));
 sky130_fd_sc_hd__o21a_1 _08807_ (.A1(net427),
    .A2(_04994_),
    .B1(_04995_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04996_));
 sky130_fd_sc_hd__mux2_1 _08808_ (.A0(\top.path[42] ),
    .A1(\top.path[43] ),
    .S(net511),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04997_));
 sky130_fd_sc_hd__o221a_1 _08809_ (.A1(\top.path[41] ),
    .A2(net325),
    .B1(_04997_),
    .B2(net426),
    .C1(net430),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04998_));
 sky130_fd_sc_hd__o21a_1 _08810_ (.A1(\top.path[40] ),
    .A2(net405),
    .B1(_04998_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_04999_));
 sky130_fd_sc_hd__mux4_1 _08811_ (.A0(\top.path[36] ),
    .A1(\top.path[37] ),
    .A2(\top.path[38] ),
    .A3(\top.path[39] ),
    .S0(net512),
    .S1(net507),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05000_));
 sky130_fd_sc_hd__mux2_1 _08812_ (.A0(\top.path[34] ),
    .A1(\top.path[35] ),
    .S(net510),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05001_));
 sky130_fd_sc_hd__or2_1 _08813_ (.A(net426),
    .B(_05001_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05002_));
 sky130_fd_sc_hd__o221a_1 _08814_ (.A1(\top.path[32] ),
    .A2(net405),
    .B1(net325),
    .B2(\top.path[33] ),
    .C1(net430),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05003_));
 sky130_fd_sc_hd__mux4_1 _08815_ (.A0(\top.path[108] ),
    .A1(\top.path[109] ),
    .A2(\top.path[110] ),
    .A3(\top.path[111] ),
    .S0(net511),
    .S1(net507),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05004_));
 sky130_fd_sc_hd__mux2_1 _08816_ (.A0(\top.path[106] ),
    .A1(\top.path[107] ),
    .S(net510),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05005_));
 sky130_fd_sc_hd__o221a_1 _08817_ (.A1(\top.path[104] ),
    .A2(net405),
    .B1(net325),
    .B2(\top.path[105] ),
    .C1(net430),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05006_));
 sky130_fd_sc_hd__o21a_1 _08818_ (.A1(net427),
    .A2(_05005_),
    .B1(_05006_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05007_));
 sky130_fd_sc_hd__a21oi_1 _08819_ (.A1(net505),
    .A2(_05004_),
    .B1(_05007_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05008_));
 sky130_fd_sc_hd__mux2_1 _08820_ (.A0(\top.path[102] ),
    .A1(\top.path[103] ),
    .S(net512),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05009_));
 sky130_fd_sc_hd__o221a_1 _08821_ (.A1(\top.path[100] ),
    .A2(net405),
    .B1(net325),
    .B2(\top.path[101] ),
    .C1(net505),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05010_));
 sky130_fd_sc_hd__o21a_1 _08822_ (.A1(net427),
    .A2(_05009_),
    .B1(_05010_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05011_));
 sky130_fd_sc_hd__mux2_1 _08823_ (.A0(\top.path[98] ),
    .A1(\top.path[99] ),
    .S(net510),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05012_));
 sky130_fd_sc_hd__o221a_1 _08824_ (.A1(\top.path[97] ),
    .A2(net325),
    .B1(_05012_),
    .B2(net427),
    .C1(net430),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05013_));
 sky130_fd_sc_hd__o21a_1 _08825_ (.A1(\top.path[96] ),
    .A2(net404),
    .B1(_05013_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05014_));
 sky130_fd_sc_hd__a221o_1 _08826_ (.A1(net505),
    .A2(_05000_),
    .B1(_05002_),
    .B2(_05003_),
    .C1(net503),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05015_));
 sky130_fd_sc_hd__o31a_1 _08827_ (.A1(_02547_),
    .A2(_04996_),
    .A3(_04999_),
    .B1(\top.translation.index[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05016_));
 sky130_fd_sc_hd__a221o_1 _08828_ (.A1(_02546_),
    .A2(_04982_),
    .B1(_05015_),
    .B2(_05016_),
    .C1(\top.translation.index[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05017_));
 sky130_fd_sc_hd__o31a_1 _08829_ (.A1(net503),
    .A2(_05011_),
    .A3(_05014_),
    .B1(\top.translation.index[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05018_));
 sky130_fd_sc_hd__a21bo_1 _08830_ (.A1(net503),
    .A2(_05008_),
    .B1_N(_05018_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05019_));
 sky130_fd_sc_hd__o311ai_1 _08831_ (.A1(net430),
    .A2(_04985_),
    .A3(_04988_),
    .B1(_04993_),
    .C1(_02546_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05020_));
 sky130_fd_sc_hd__a31o_1 _08832_ (.A1(\top.translation.index[6] ),
    .A2(_05019_),
    .A3(_05020_),
    .B1(\top.translation.index[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05021_));
 sky130_fd_sc_hd__inv_2 _08833_ (.A(_05021_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05022_));
 sky130_fd_sc_hd__a32o_1 _08834_ (.A1(\top.translation.index[4] ),
    .A2(_04962_),
    .A3(_04969_),
    .B1(_05017_),
    .B2(_05022_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05023_));
 sky130_fd_sc_hd__and2b_1 _08835_ (.A_N(\top.translation.write_fin ),
    .B(\top.TRN_sram_complete ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05024_));
 sky130_fd_sc_hd__inv_2 _08836_ (.A(_05024_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05025_));
 sky130_fd_sc_hd__or4_1 _08837_ (.A(\top.TRN_char_index[6] ),
    .B(\top.TRN_char_index[5] ),
    .C(\top.TRN_char_index[0] ),
    .D(\top.TRN_sram_complete ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05026_));
 sky130_fd_sc_hd__and4b_1 _08838_ (.A_N(\top.TRN_char_index[2] ),
    .B(\top.TRN_char_index[1] ),
    .C(\top.TRN_char_index[4] ),
    .D(\top.TRN_char_index[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05027_));
 sky130_fd_sc_hd__and2b_1 _08839_ (.A_N(_05026_),
    .B(_05027_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05028_));
 sky130_fd_sc_hd__or4_1 _08840_ (.A(net513),
    .B(\top.translation.totalEn ),
    .C(net466),
    .D(_05028_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05029_));
 sky130_fd_sc_hd__or4_1 _08841_ (.A(_02813_),
    .B(_05023_),
    .C(_05025_),
    .D(_05029_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05030_));
 sky130_fd_sc_hd__o211a_1 _08842_ (.A1(net423),
    .A2(\top.header_synthesis.enable ),
    .B1(net36),
    .C1(net452),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05031_));
 sky130_fd_sc_hd__o211a_1 _08843_ (.A1(_05024_),
    .A2(_05029_),
    .B1(_05030_),
    .C1(_05031_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05032_));
 sky130_fd_sc_hd__o21ba_1 _08844_ (.A1(_02813_),
    .A2(_05028_),
    .B1_N(\top.translation.totalEn ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05033_));
 sky130_fd_sc_hd__o21ai_1 _08845_ (.A1(net513),
    .A2(_05033_),
    .B1(net423),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05034_));
 sky130_fd_sc_hd__mux2_1 _08846_ (.A0(net1103),
    .A1(_05034_),
    .S(_05032_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01449_));
 sky130_fd_sc_hd__or3_1 _08847_ (.A(net513),
    .B(\top.translation.totalEn ),
    .C(_05024_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05035_));
 sky130_fd_sc_hd__and3_1 _08848_ (.A(net452),
    .B(_02807_),
    .C(_05035_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05036_));
 sky130_fd_sc_hd__nand2_1 _08849_ (.A(_02808_),
    .B(_05035_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05037_));
 sky130_fd_sc_hd__o21a_1 _08850_ (.A1(\top.translation.index[5] ),
    .A2(_02812_),
    .B1(\top.translation.index[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05038_));
 sky130_fd_sc_hd__nand2_1 _08851_ (.A(_02550_),
    .B(_05036_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05039_));
 sky130_fd_sc_hd__o32a_1 _08852_ (.A1(_02813_),
    .A2(_05038_),
    .A3(_05039_),
    .B1(_05036_),
    .B2(\top.translation.index[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01448_));
 sky130_fd_sc_hd__a21oi_1 _08853_ (.A1(_02550_),
    .A2(_02812_),
    .B1(_05037_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05040_));
 sky130_fd_sc_hd__or2_1 _08854_ (.A(\top.translation.index[5] ),
    .B(_05040_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05041_));
 sky130_fd_sc_hd__o31a_1 _08855_ (.A1(_02546_),
    .A2(_02812_),
    .A3(_05039_),
    .B1(_05041_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01447_));
 sky130_fd_sc_hd__or3b_1 _08856_ (.A(_05037_),
    .B(net502),
    .C_N(_02811_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05042_));
 sky130_fd_sc_hd__a21o_1 _08857_ (.A1(\top.translation.index[4] ),
    .A2(_05042_),
    .B1(_05040_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01446_));
 sky130_fd_sc_hd__o21a_1 _08858_ (.A1(net513),
    .A2(_02811_),
    .B1(_05036_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05043_));
 sky130_fd_sc_hd__nand2_1 _08859_ (.A(net502),
    .B(_02811_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05044_));
 sky130_fd_sc_hd__o22a_1 _08860_ (.A1(net502),
    .A2(_05043_),
    .B1(_05044_),
    .B2(_05039_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01445_));
 sky130_fd_sc_hd__o21a_1 _08861_ (.A1(net402),
    .A2(_05037_),
    .B1(net504),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05045_));
 sky130_fd_sc_hd__or2_1 _08862_ (.A(_05043_),
    .B(_05045_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01444_));
 sky130_fd_sc_hd__or2_1 _08863_ (.A(net509),
    .B(_05037_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05046_));
 sky130_fd_sc_hd__and2_1 _08864_ (.A(_02550_),
    .B(net402),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05047_));
 sky130_fd_sc_hd__a2bb2o_1 _08865_ (.A1_N(_05047_),
    .A2_N(_05037_),
    .B1(net506),
    .B2(_05046_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01443_));
 sky130_fd_sc_hd__a21bo_1 _08866_ (.A1(net509),
    .A2(_05039_),
    .B1_N(_05046_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01442_));
 sky130_fd_sc_hd__a21o_1 _08867_ (.A1(_02808_),
    .A2(_02813_),
    .B1(net513),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05048_));
 sky130_fd_sc_hd__nand2_1 _08868_ (.A(net513),
    .B(_02808_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05049_));
 sky130_fd_sc_hd__and3_1 _08869_ (.A(_05035_),
    .B(_05048_),
    .C(_05049_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01441_));
 sky130_fd_sc_hd__and2_1 _08870_ (.A(\top.translation.totalEn ),
    .B(_05049_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01440_));
 sky130_fd_sc_hd__mux2_1 _08871_ (.A0(net1057),
    .A1(\top.WB.CPU_DAT_O[31] ),
    .S(net303),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01439_));
 sky130_fd_sc_hd__mux2_1 _08872_ (.A0(net1062),
    .A1(\top.WB.CPU_DAT_O[30] ),
    .S(net303),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01438_));
 sky130_fd_sc_hd__mux2_1 _08873_ (.A0(net1116),
    .A1(\top.WB.CPU_DAT_O[29] ),
    .S(net303),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01437_));
 sky130_fd_sc_hd__mux2_1 _08874_ (.A0(net1156),
    .A1(\top.WB.CPU_DAT_O[28] ),
    .S(net303),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01436_));
 sky130_fd_sc_hd__mux2_1 _08875_ (.A0(net1114),
    .A1(\top.WB.CPU_DAT_O[27] ),
    .S(net302),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01435_));
 sky130_fd_sc_hd__mux2_1 _08876_ (.A0(net1060),
    .A1(\top.WB.CPU_DAT_O[26] ),
    .S(net302),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01434_));
 sky130_fd_sc_hd__mux2_1 _08877_ (.A0(net1337),
    .A1(\top.WB.CPU_DAT_O[25] ),
    .S(net302),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01433_));
 sky130_fd_sc_hd__mux2_1 _08878_ (.A0(net1190),
    .A1(\top.WB.CPU_DAT_O[24] ),
    .S(net302),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01432_));
 sky130_fd_sc_hd__mux2_1 _08879_ (.A0(net1055),
    .A1(\top.WB.CPU_DAT_O[23] ),
    .S(net303),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01431_));
 sky130_fd_sc_hd__mux2_1 _08880_ (.A0(net1046),
    .A1(\top.WB.CPU_DAT_O[22] ),
    .S(net303),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01430_));
 sky130_fd_sc_hd__mux2_1 _08881_ (.A0(net1326),
    .A1(\top.WB.CPU_DAT_O[21] ),
    .S(net302),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01429_));
 sky130_fd_sc_hd__mux2_1 _08882_ (.A0(net1207),
    .A1(\top.WB.CPU_DAT_O[20] ),
    .S(net302),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01428_));
 sky130_fd_sc_hd__mux2_1 _08883_ (.A0(net1106),
    .A1(\top.WB.CPU_DAT_O[19] ),
    .S(net302),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01427_));
 sky130_fd_sc_hd__mux2_1 _08884_ (.A0(net1069),
    .A1(\top.WB.CPU_DAT_O[18] ),
    .S(net302),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01426_));
 sky130_fd_sc_hd__mux2_1 _08885_ (.A0(net1442),
    .A1(\top.WB.CPU_DAT_O[17] ),
    .S(net302),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01425_));
 sky130_fd_sc_hd__mux2_1 _08886_ (.A0(net1162),
    .A1(\top.WB.CPU_DAT_O[16] ),
    .S(net302),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01424_));
 sky130_fd_sc_hd__mux2_1 _08887_ (.A0(net1200),
    .A1(\top.WB.CPU_DAT_O[15] ),
    .S(net305),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01423_));
 sky130_fd_sc_hd__mux2_1 _08888_ (.A0(net1218),
    .A1(\top.WB.CPU_DAT_O[14] ),
    .S(net305),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01422_));
 sky130_fd_sc_hd__mux2_1 _08889_ (.A0(net1407),
    .A1(\top.WB.CPU_DAT_O[13] ),
    .S(net306),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01421_));
 sky130_fd_sc_hd__mux2_1 _08890_ (.A0(net1224),
    .A1(\top.WB.CPU_DAT_O[12] ),
    .S(net306),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01420_));
 sky130_fd_sc_hd__mux2_1 _08891_ (.A0(net1159),
    .A1(\top.WB.CPU_DAT_O[11] ),
    .S(net305),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01419_));
 sky130_fd_sc_hd__mux2_1 _08892_ (.A0(net1084),
    .A1(\top.WB.CPU_DAT_O[10] ),
    .S(net306),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01418_));
 sky130_fd_sc_hd__mux2_1 _08893_ (.A0(net1308),
    .A1(\top.WB.CPU_DAT_O[9] ),
    .S(net305),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01417_));
 sky130_fd_sc_hd__mux2_1 _08894_ (.A0(net1044),
    .A1(\top.WB.CPU_DAT_O[8] ),
    .S(net306),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01416_));
 sky130_fd_sc_hd__mux2_1 _08895_ (.A0(net1078),
    .A1(\top.WB.CPU_DAT_O[7] ),
    .S(net305),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01415_));
 sky130_fd_sc_hd__mux2_1 _08896_ (.A0(net1091),
    .A1(\top.WB.CPU_DAT_O[6] ),
    .S(net305),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01414_));
 sky130_fd_sc_hd__mux2_1 _08897_ (.A0(net1110),
    .A1(\top.WB.CPU_DAT_O[5] ),
    .S(net305),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01413_));
 sky130_fd_sc_hd__mux2_1 _08898_ (.A0(net1148),
    .A1(\top.WB.CPU_DAT_O[4] ),
    .S(net306),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01412_));
 sky130_fd_sc_hd__mux2_1 _08899_ (.A0(net1054),
    .A1(\top.WB.CPU_DAT_O[3] ),
    .S(net305),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01411_));
 sky130_fd_sc_hd__mux2_1 _08900_ (.A0(net1187),
    .A1(\top.WB.CPU_DAT_O[2] ),
    .S(net305),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01410_));
 sky130_fd_sc_hd__mux2_1 _08901_ (.A0(net1240),
    .A1(\top.WB.CPU_DAT_O[1] ),
    .S(net306),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01409_));
 sky130_fd_sc_hd__mux2_1 _08902_ (.A0(net1239),
    .A1(\top.WB.CPU_DAT_O[0] ),
    .S(net305),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01408_));
 sky130_fd_sc_hd__or2_1 _08903_ (.A(_02522_),
    .B(_02831_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05050_));
 sky130_fd_sc_hd__nor3_1 _08904_ (.A(_02418_),
    .B(net422),
    .C(_05050_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05051_));
 sky130_fd_sc_hd__nor2_1 _08905_ (.A(net470),
    .B(_02851_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05052_));
 sky130_fd_sc_hd__a311o_1 _08906_ (.A1(_02418_),
    .A2(\top.hTree.closing ),
    .A3(net470),
    .B1(_05051_),
    .C1(_05052_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05053_));
 sky130_fd_sc_hd__nand2_1 _08907_ (.A(net288),
    .B(_04255_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05054_));
 sky130_fd_sc_hd__o2bb2a_1 _08908_ (.A1_N(\top.hTree.finish_check ),
    .A2_N(_04254_),
    .B1(_05053_),
    .B2(_05054_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05055_));
 sky130_fd_sc_hd__and3b_1 _08909_ (.A_N(_02835_),
    .B(_05050_),
    .C(\top.findLeastValue.least2[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05056_));
 sky130_fd_sc_hd__and3_1 _08910_ (.A(\top.hTree.write_HT_fin ),
    .B(net470),
    .C(_05056_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05057_));
 sky130_fd_sc_hd__nand2_1 _08911_ (.A(net449),
    .B(_02838_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05058_));
 sky130_fd_sc_hd__or4_4 _08912_ (.A(_02866_),
    .B(_05055_),
    .C(_05057_),
    .D(_05058_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05059_));
 sky130_fd_sc_hd__and4_1 _08913_ (.A(\top.cb_syn.max_index[4] ),
    .B(\top.cb_syn.max_index[3] ),
    .C(\top.cb_syn.max_index[2] ),
    .D(\top.cb_syn.max_index[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05060_));
 sky130_fd_sc_hd__and3_1 _08914_ (.A(\top.cb_syn.max_index[6] ),
    .B(\top.cb_syn.max_index[5] ),
    .C(_05060_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05061_));
 sky130_fd_sc_hd__xor2_1 _08915_ (.A(\top.cb_syn.max_index[7] ),
    .B(_05061_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05062_));
 sky130_fd_sc_hd__mux2_1 _08916_ (.A0(_04186_),
    .A1(_05062_),
    .S(_04255_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05063_));
 sky130_fd_sc_hd__mux2_1 _08917_ (.A0(_05063_),
    .A1(\top.cb_syn.max_index[7] ),
    .S(_05059_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01407_));
 sky130_fd_sc_hd__a21oi_1 _08918_ (.A1(\top.cb_syn.max_index[5] ),
    .A2(_05060_),
    .B1(\top.cb_syn.max_index[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05064_));
 sky130_fd_sc_hd__nor2_1 _08919_ (.A(_05061_),
    .B(_05064_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05065_));
 sky130_fd_sc_hd__mux2_1 _08920_ (.A0(_04217_),
    .A1(_05065_),
    .S(_04255_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05066_));
 sky130_fd_sc_hd__mux2_1 _08921_ (.A0(_05066_),
    .A1(\top.cb_syn.max_index[6] ),
    .S(_05059_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01406_));
 sky130_fd_sc_hd__xor2_1 _08922_ (.A(\top.cb_syn.max_index[5] ),
    .B(_05060_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05067_));
 sky130_fd_sc_hd__mux2_1 _08923_ (.A0(_04222_),
    .A1(_05067_),
    .S(_04255_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05068_));
 sky130_fd_sc_hd__mux2_1 _08924_ (.A0(_05068_),
    .A1(\top.cb_syn.max_index[5] ),
    .S(_05059_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01405_));
 sky130_fd_sc_hd__a31o_1 _08925_ (.A1(\top.cb_syn.max_index[3] ),
    .A2(\top.cb_syn.max_index[2] ),
    .A3(\top.cb_syn.max_index[1] ),
    .B1(\top.cb_syn.max_index[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05069_));
 sky130_fd_sc_hd__or3b_1 _08926_ (.A(_04254_),
    .B(_05060_),
    .C_N(_05069_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05070_));
 sky130_fd_sc_hd__a21bo_1 _08927_ (.A1(_04228_),
    .A2(_04254_),
    .B1_N(_05070_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05071_));
 sky130_fd_sc_hd__mux2_1 _08928_ (.A0(_05071_),
    .A1(\top.cb_syn.max_index[4] ),
    .S(_05059_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01404_));
 sky130_fd_sc_hd__nand2_1 _08929_ (.A(_04240_),
    .B(_04255_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05072_));
 sky130_fd_sc_hd__xnor2_1 _08930_ (.A(_04234_),
    .B(_05072_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05073_));
 sky130_fd_sc_hd__mux2_1 _08931_ (.A0(_05073_),
    .A1(\top.cb_syn.max_index[3] ),
    .S(_05059_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01403_));
 sky130_fd_sc_hd__a21oi_1 _08932_ (.A1(_04239_),
    .A2(_04254_),
    .B1(_05059_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05074_));
 sky130_fd_sc_hd__a22o_1 _08933_ (.A1(\top.cb_syn.max_index[2] ),
    .A2(_05059_),
    .B1(_05072_),
    .B2(_05074_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01402_));
 sky130_fd_sc_hd__xnor2_1 _08934_ (.A(\top.cb_syn.max_index[1] ),
    .B(_05059_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_01401_));
 sky130_fd_sc_hd__or4b_2 _08935_ (.A(\top.sram_interface.TRN_counter[2] ),
    .B(\top.sram_interface.TRN_counter[0] ),
    .C(_02914_),
    .D_N(\top.sram_interface.TRN_counter[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05075_));
 sky130_fd_sc_hd__inv_2 _08936_ (.A(_05075_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05076_));
 sky130_fd_sc_hd__mux2_1 _08937_ (.A0(\top.WB.CPU_DAT_O[31] ),
    .A1(net1393),
    .S(net319),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01400_));
 sky130_fd_sc_hd__mux2_1 _08938_ (.A0(\top.WB.CPU_DAT_O[30] ),
    .A1(net1289),
    .S(net319),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01399_));
 sky130_fd_sc_hd__mux2_1 _08939_ (.A0(\top.WB.CPU_DAT_O[29] ),
    .A1(net1414),
    .S(net319),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01398_));
 sky130_fd_sc_hd__mux2_1 _08940_ (.A0(\top.WB.CPU_DAT_O[28] ),
    .A1(net1468),
    .S(net318),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01397_));
 sky130_fd_sc_hd__mux2_1 _08941_ (.A0(\top.WB.CPU_DAT_O[27] ),
    .A1(net1267),
    .S(net319),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01396_));
 sky130_fd_sc_hd__mux2_1 _08942_ (.A0(\top.WB.CPU_DAT_O[26] ),
    .A1(net1265),
    .S(net318),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01395_));
 sky130_fd_sc_hd__mux2_1 _08943_ (.A0(\top.WB.CPU_DAT_O[25] ),
    .A1(net1374),
    .S(net322),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01394_));
 sky130_fd_sc_hd__mux2_1 _08944_ (.A0(\top.WB.CPU_DAT_O[24] ),
    .A1(net1389),
    .S(net322),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01393_));
 sky130_fd_sc_hd__mux2_1 _08945_ (.A0(\top.WB.CPU_DAT_O[23] ),
    .A1(net1254),
    .S(net318),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01392_));
 sky130_fd_sc_hd__mux2_1 _08946_ (.A0(\top.WB.CPU_DAT_O[22] ),
    .A1(net1215),
    .S(net318),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01391_));
 sky130_fd_sc_hd__mux2_1 _08947_ (.A0(\top.WB.CPU_DAT_O[21] ),
    .A1(net1419),
    .S(net318),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01390_));
 sky130_fd_sc_hd__mux2_1 _08948_ (.A0(\top.WB.CPU_DAT_O[20] ),
    .A1(net1435),
    .S(net318),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01389_));
 sky130_fd_sc_hd__mux2_1 _08949_ (.A0(\top.WB.CPU_DAT_O[19] ),
    .A1(net1124),
    .S(net318),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01388_));
 sky130_fd_sc_hd__mux2_1 _08950_ (.A0(\top.WB.CPU_DAT_O[18] ),
    .A1(net1165),
    .S(net318),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01387_));
 sky130_fd_sc_hd__mux2_1 _08951_ (.A0(\top.WB.CPU_DAT_O[17] ),
    .A1(net1065),
    .S(net318),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01386_));
 sky130_fd_sc_hd__mux2_1 _08952_ (.A0(\top.WB.CPU_DAT_O[16] ),
    .A1(net1341),
    .S(net318),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01385_));
 sky130_fd_sc_hd__mux2_1 _08953_ (.A0(\top.WB.CPU_DAT_O[15] ),
    .A1(net1381),
    .S(net321),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01384_));
 sky130_fd_sc_hd__mux2_1 _08954_ (.A0(\top.WB.CPU_DAT_O[14] ),
    .A1(net1398),
    .S(net321),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01383_));
 sky130_fd_sc_hd__mux2_1 _08955_ (.A0(\top.WB.CPU_DAT_O[13] ),
    .A1(net1253),
    .S(net320),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01382_));
 sky130_fd_sc_hd__mux2_1 _08956_ (.A0(\top.WB.CPU_DAT_O[12] ),
    .A1(net1217),
    .S(net320),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01381_));
 sky130_fd_sc_hd__mux2_1 _08957_ (.A0(\top.WB.CPU_DAT_O[11] ),
    .A1(net1345),
    .S(net320),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01380_));
 sky130_fd_sc_hd__mux2_1 _08958_ (.A0(\top.WB.CPU_DAT_O[10] ),
    .A1(net1394),
    .S(net320),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01379_));
 sky130_fd_sc_hd__mux2_1 _08959_ (.A0(\top.WB.CPU_DAT_O[9] ),
    .A1(net1453),
    .S(net320),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01378_));
 sky130_fd_sc_hd__mux2_1 _08960_ (.A0(\top.WB.CPU_DAT_O[8] ),
    .A1(net1146),
    .S(net320),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01377_));
 sky130_fd_sc_hd__mux2_1 _08961_ (.A0(\top.WB.CPU_DAT_O[7] ),
    .A1(net1234),
    .S(net321),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01376_));
 sky130_fd_sc_hd__mux2_1 _08962_ (.A0(\top.WB.CPU_DAT_O[6] ),
    .A1(net1257),
    .S(net321),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01375_));
 sky130_fd_sc_hd__mux2_1 _08963_ (.A0(\top.WB.CPU_DAT_O[5] ),
    .A1(net1380),
    .S(net321),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01374_));
 sky130_fd_sc_hd__mux2_1 _08964_ (.A0(\top.WB.CPU_DAT_O[4] ),
    .A1(net1352),
    .S(net321),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01373_));
 sky130_fd_sc_hd__mux2_1 _08965_ (.A0(\top.WB.CPU_DAT_O[3] ),
    .A1(net1250),
    .S(net320),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01372_));
 sky130_fd_sc_hd__mux2_1 _08966_ (.A0(\top.WB.CPU_DAT_O[2] ),
    .A1(net1258),
    .S(net320),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01371_));
 sky130_fd_sc_hd__mux2_1 _08967_ (.A0(\top.WB.CPU_DAT_O[1] ),
    .A1(net1377),
    .S(net320),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01370_));
 sky130_fd_sc_hd__mux2_1 _08968_ (.A0(\top.WB.CPU_DAT_O[0] ),
    .A1(net1401),
    .S(net320),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01369_));
 sky130_fd_sc_hd__nand2_1 _08969_ (.A(net465),
    .B(\top.sram_interface.word_cnt[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05077_));
 sky130_fd_sc_hd__mux2_1 _08970_ (.A0(\top.WB.CPU_DAT_O[31] ),
    .A1(net550),
    .S(net368),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01368_));
 sky130_fd_sc_hd__mux2_1 _08971_ (.A0(\top.WB.CPU_DAT_O[30] ),
    .A1(net1598),
    .S(net368),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01367_));
 sky130_fd_sc_hd__mux2_1 _08972_ (.A0(\top.WB.CPU_DAT_O[29] ),
    .A1(\top.cb_syn.h_element[61] ),
    .S(net367),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01366_));
 sky130_fd_sc_hd__mux2_1 _08973_ (.A0(\top.WB.CPU_DAT_O[28] ),
    .A1(\top.cb_syn.h_element[60] ),
    .S(net368),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01365_));
 sky130_fd_sc_hd__mux2_1 _08974_ (.A0(\top.WB.CPU_DAT_O[27] ),
    .A1(\top.cb_syn.h_element[59] ),
    .S(net367),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01364_));
 sky130_fd_sc_hd__mux2_1 _08975_ (.A0(\top.WB.CPU_DAT_O[26] ),
    .A1(net1769),
    .S(net367),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01363_));
 sky130_fd_sc_hd__mux2_1 _08976_ (.A0(\top.WB.CPU_DAT_O[25] ),
    .A1(\top.cb_syn.h_element[57] ),
    .S(net367),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01362_));
 sky130_fd_sc_hd__mux2_1 _08977_ (.A0(\top.WB.CPU_DAT_O[24] ),
    .A1(net1780),
    .S(net367),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01361_));
 sky130_fd_sc_hd__mux2_1 _08978_ (.A0(\top.WB.CPU_DAT_O[23] ),
    .A1(\top.cb_syn.h_element[55] ),
    .S(net368),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01360_));
 sky130_fd_sc_hd__mux2_1 _08979_ (.A0(\top.WB.CPU_DAT_O[22] ),
    .A1(\top.cb_syn.h_element[54] ),
    .S(net368),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01359_));
 sky130_fd_sc_hd__mux2_1 _08980_ (.A0(\top.WB.CPU_DAT_O[21] ),
    .A1(net1485),
    .S(net367),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01358_));
 sky130_fd_sc_hd__mux2_1 _08981_ (.A0(\top.WB.CPU_DAT_O[20] ),
    .A1(\top.cb_syn.h_element[52] ),
    .S(net368),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01357_));
 sky130_fd_sc_hd__mux2_1 _08982_ (.A0(\top.WB.CPU_DAT_O[19] ),
    .A1(\top.cb_syn.h_element[51] ),
    .S(net367),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01356_));
 sky130_fd_sc_hd__mux2_1 _08983_ (.A0(\top.WB.CPU_DAT_O[18] ),
    .A1(\top.cb_syn.h_element[50] ),
    .S(net367),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01355_));
 sky130_fd_sc_hd__mux2_1 _08984_ (.A0(\top.WB.CPU_DAT_O[17] ),
    .A1(\top.cb_syn.h_element[49] ),
    .S(net367),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01354_));
 sky130_fd_sc_hd__mux2_1 _08985_ (.A0(\top.WB.CPU_DAT_O[16] ),
    .A1(\top.cb_syn.h_element[48] ),
    .S(net367),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01353_));
 sky130_fd_sc_hd__mux2_1 _08986_ (.A0(\top.WB.CPU_DAT_O[15] ),
    .A1(\top.cb_syn.h_element[47] ),
    .S(net368),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01352_));
 sky130_fd_sc_hd__mux2_1 _08987_ (.A0(\top.WB.CPU_DAT_O[14] ),
    .A1(\top.cb_syn.h_element[46] ),
    .S(net368),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01351_));
 sky130_fd_sc_hd__nand2_1 _08988_ (.A(net449),
    .B(net528),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05078_));
 sky130_fd_sc_hd__mux2_1 _08989_ (.A0(\top.WB.CPU_DAT_O[31] ),
    .A1(net1301),
    .S(net366),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01350_));
 sky130_fd_sc_hd__mux2_1 _08990_ (.A0(\top.WB.CPU_DAT_O[30] ),
    .A1(net1206),
    .S(net366),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01349_));
 sky130_fd_sc_hd__mux2_1 _08991_ (.A0(\top.WB.CPU_DAT_O[29] ),
    .A1(net1268),
    .S(net366),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01348_));
 sky130_fd_sc_hd__mux2_1 _08992_ (.A0(\top.WB.CPU_DAT_O[28] ),
    .A1(net1249),
    .S(net366),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01347_));
 sky130_fd_sc_hd__mux2_1 _08993_ (.A0(\top.WB.CPU_DAT_O[27] ),
    .A1(net1164),
    .S(net366),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01346_));
 sky130_fd_sc_hd__mux2_1 _08994_ (.A0(\top.WB.CPU_DAT_O[26] ),
    .A1(net1192),
    .S(net365),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01345_));
 sky130_fd_sc_hd__mux2_1 _08995_ (.A0(\top.WB.CPU_DAT_O[25] ),
    .A1(net1344),
    .S(net365),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01344_));
 sky130_fd_sc_hd__mux2_1 _08996_ (.A0(\top.WB.CPU_DAT_O[24] ),
    .A1(net1340),
    .S(net366),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01343_));
 sky130_fd_sc_hd__mux2_1 _08997_ (.A0(\top.WB.CPU_DAT_O[23] ),
    .A1(net1335),
    .S(net365),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01342_));
 sky130_fd_sc_hd__mux2_1 _08998_ (.A0(\top.WB.CPU_DAT_O[22] ),
    .A1(net1212),
    .S(net366),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01341_));
 sky130_fd_sc_hd__mux2_1 _08999_ (.A0(\top.WB.CPU_DAT_O[21] ),
    .A1(net1168),
    .S(net365),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01340_));
 sky130_fd_sc_hd__mux2_1 _09000_ (.A0(\top.WB.CPU_DAT_O[20] ),
    .A1(net1425),
    .S(net365),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01339_));
 sky130_fd_sc_hd__mux2_1 _09001_ (.A0(\top.WB.CPU_DAT_O[19] ),
    .A1(net1486),
    .S(net365),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01338_));
 sky130_fd_sc_hd__mux2_1 _09002_ (.A0(\top.WB.CPU_DAT_O[18] ),
    .A1(net1445),
    .S(net365),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01337_));
 sky130_fd_sc_hd__mux2_1 _09003_ (.A0(\top.WB.CPU_DAT_O[17] ),
    .A1(net1260),
    .S(net365),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01336_));
 sky130_fd_sc_hd__mux2_1 _09004_ (.A0(\top.WB.CPU_DAT_O[16] ),
    .A1(net1222),
    .S(net365),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01335_));
 sky130_fd_sc_hd__mux2_1 _09005_ (.A0(\top.WB.CPU_DAT_O[15] ),
    .A1(net1331),
    .S(net366),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01334_));
 sky130_fd_sc_hd__mux2_1 _09006_ (.A0(\top.WB.CPU_DAT_O[14] ),
    .A1(net1270),
    .S(net365),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01333_));
 sky130_fd_sc_hd__and2_1 _09007_ (.A(\top.histogram.eof_n ),
    .B(_03321_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05079_));
 sky130_fd_sc_hd__nor2_2 _09008_ (.A(net444),
    .B(_02405_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05080_));
 sky130_fd_sc_hd__o31ai_4 _09009_ (.A1(_03364_),
    .A2(_05079_),
    .A3(_05080_),
    .B1(net453),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05081_));
 sky130_fd_sc_hd__o21ba_2 _09010_ (.A1(\top.histogram.eof_n ),
    .A2(_05080_),
    .B1_N(_05081_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05082_));
 sky130_fd_sc_hd__a22o_1 _09011_ (.A1(net1685),
    .A2(_05081_),
    .B1(_05082_),
    .B2(\top.TRN_char_index[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01332_));
 sky130_fd_sc_hd__a22o_1 _09012_ (.A1(net1575),
    .A2(_05081_),
    .B1(_05082_),
    .B2(\top.TRN_char_index[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01331_));
 sky130_fd_sc_hd__a22o_1 _09013_ (.A1(net1758),
    .A2(_05081_),
    .B1(_05082_),
    .B2(\top.TRN_char_index[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01330_));
 sky130_fd_sc_hd__a22o_1 _09014_ (.A1(net1612),
    .A2(_05081_),
    .B1(_05082_),
    .B2(\top.TRN_char_index[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01329_));
 sky130_fd_sc_hd__a22o_1 _09015_ (.A1(\top.hist_addr[2] ),
    .A2(_05081_),
    .B1(_05082_),
    .B2(net445),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01328_));
 sky130_fd_sc_hd__a22o_1 _09016_ (.A1(net1797),
    .A2(_05081_),
    .B1(_05082_),
    .B2(\top.TRN_char_index[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01327_));
 sky130_fd_sc_hd__a22o_1 _09017_ (.A1(net1740),
    .A2(_05081_),
    .B1(_05082_),
    .B2(\top.TRN_char_index[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01326_));
 sky130_fd_sc_hd__or4b_1 _09018_ (.A(\top.sram_interface.TRN_counter[2] ),
    .B(_02914_),
    .C(\top.sram_interface.TRN_counter[1] ),
    .D_N(\top.sram_interface.TRN_counter[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05083_));
 sky130_fd_sc_hd__mux2_1 _09019_ (.A0(\top.WB.CPU_DAT_O[31] ),
    .A1(net1306),
    .S(net314),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01325_));
 sky130_fd_sc_hd__mux2_1 _09020_ (.A0(\top.WB.CPU_DAT_O[30] ),
    .A1(net1135),
    .S(net314),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01324_));
 sky130_fd_sc_hd__mux2_1 _09021_ (.A0(\top.WB.CPU_DAT_O[29] ),
    .A1(net1328),
    .S(net314),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01323_));
 sky130_fd_sc_hd__mux2_1 _09022_ (.A0(\top.WB.CPU_DAT_O[28] ),
    .A1(net1372),
    .S(net313),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01322_));
 sky130_fd_sc_hd__mux2_1 _09023_ (.A0(\top.WB.CPU_DAT_O[27] ),
    .A1(net1223),
    .S(net314),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01321_));
 sky130_fd_sc_hd__mux2_1 _09024_ (.A0(\top.WB.CPU_DAT_O[26] ),
    .A1(net1279),
    .S(net314),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01320_));
 sky130_fd_sc_hd__mux2_1 _09025_ (.A0(\top.WB.CPU_DAT_O[25] ),
    .A1(net1194),
    .S(net313),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01319_));
 sky130_fd_sc_hd__mux2_1 _09026_ (.A0(\top.WB.CPU_DAT_O[24] ),
    .A1(net1294),
    .S(net313),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01318_));
 sky130_fd_sc_hd__mux2_1 _09027_ (.A0(\top.WB.CPU_DAT_O[23] ),
    .A1(net1205),
    .S(net313),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01317_));
 sky130_fd_sc_hd__mux2_1 _09028_ (.A0(\top.WB.CPU_DAT_O[22] ),
    .A1(net1107),
    .S(net314),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01316_));
 sky130_fd_sc_hd__mux2_1 _09029_ (.A0(\top.WB.CPU_DAT_O[21] ),
    .A1(net1403),
    .S(net313),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01315_));
 sky130_fd_sc_hd__mux2_1 _09030_ (.A0(\top.WB.CPU_DAT_O[20] ),
    .A1(net1382),
    .S(net313),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01314_));
 sky130_fd_sc_hd__mux2_1 _09031_ (.A0(\top.WB.CPU_DAT_O[19] ),
    .A1(net1202),
    .S(net313),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01313_));
 sky130_fd_sc_hd__mux2_1 _09032_ (.A0(\top.WB.CPU_DAT_O[18] ),
    .A1(net1300),
    .S(net313),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01312_));
 sky130_fd_sc_hd__mux2_1 _09033_ (.A0(\top.WB.CPU_DAT_O[17] ),
    .A1(net1263),
    .S(net313),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01311_));
 sky130_fd_sc_hd__mux2_1 _09034_ (.A0(\top.WB.CPU_DAT_O[16] ),
    .A1(net1144),
    .S(net313),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01310_));
 sky130_fd_sc_hd__mux2_1 _09035_ (.A0(\top.WB.CPU_DAT_O[15] ),
    .A1(net1134),
    .S(net315),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01309_));
 sky130_fd_sc_hd__mux2_1 _09036_ (.A0(\top.WB.CPU_DAT_O[14] ),
    .A1(net1286),
    .S(net315),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01308_));
 sky130_fd_sc_hd__mux2_1 _09037_ (.A0(\top.WB.CPU_DAT_O[13] ),
    .A1(net1181),
    .S(net315),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01307_));
 sky130_fd_sc_hd__mux2_1 _09038_ (.A0(\top.WB.CPU_DAT_O[12] ),
    .A1(net1095),
    .S(net315),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01306_));
 sky130_fd_sc_hd__mux2_1 _09039_ (.A0(\top.WB.CPU_DAT_O[11] ),
    .A1(net1259),
    .S(net315),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01305_));
 sky130_fd_sc_hd__mux2_1 _09040_ (.A0(\top.WB.CPU_DAT_O[10] ),
    .A1(net1311),
    .S(net315),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01304_));
 sky130_fd_sc_hd__mux2_1 _09041_ (.A0(\top.WB.CPU_DAT_O[9] ),
    .A1(net1496),
    .S(net315),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01303_));
 sky130_fd_sc_hd__mux2_1 _09042_ (.A0(\top.WB.CPU_DAT_O[8] ),
    .A1(net1459),
    .S(net315),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01302_));
 sky130_fd_sc_hd__mux2_1 _09043_ (.A0(\top.WB.CPU_DAT_O[7] ),
    .A1(net1183),
    .S(net315),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01301_));
 sky130_fd_sc_hd__mux2_1 _09044_ (.A0(\top.WB.CPU_DAT_O[6] ),
    .A1(net1315),
    .S(net316),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01300_));
 sky130_fd_sc_hd__mux2_1 _09045_ (.A0(\top.WB.CPU_DAT_O[5] ),
    .A1(net1406),
    .S(net315),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01299_));
 sky130_fd_sc_hd__mux2_1 _09046_ (.A0(\top.WB.CPU_DAT_O[4] ),
    .A1(net1369),
    .S(net316),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01298_));
 sky130_fd_sc_hd__mux2_1 _09047_ (.A0(\top.WB.CPU_DAT_O[3] ),
    .A1(net1418),
    .S(net316),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01297_));
 sky130_fd_sc_hd__mux2_1 _09048_ (.A0(\top.WB.CPU_DAT_O[2] ),
    .A1(net1373),
    .S(net316),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01296_));
 sky130_fd_sc_hd__mux2_1 _09049_ (.A0(\top.WB.CPU_DAT_O[1] ),
    .A1(net1471),
    .S(net316),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01295_));
 sky130_fd_sc_hd__mux2_1 _09050_ (.A0(\top.WB.CPU_DAT_O[0] ),
    .A1(net1533),
    .S(net316),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01294_));
 sky130_fd_sc_hd__or3_1 _09051_ (.A(_02552_),
    .B(_02882_),
    .C(_02883_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05084_));
 sky130_fd_sc_hd__nor2_1 _09052_ (.A(net412),
    .B(_05084_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05085_));
 sky130_fd_sc_hd__or2_1 _09053_ (.A(net412),
    .B(_05084_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05086_));
 sky130_fd_sc_hd__a22o_1 _09054_ (.A1(\top.cb_syn.char_path_n[1] ),
    .A2(_04202_),
    .B1(_04585_),
    .B2(_05085_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05087_));
 sky130_fd_sc_hd__a31o_1 _09055_ (.A1(\top.CB_write_complete ),
    .A2(\top.cb_syn.end_cond ),
    .A3(\top.cb_syn.curr_state[8] ),
    .B1(_05087_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05088_));
 sky130_fd_sc_hd__a21o_1 _09056_ (.A1(net463),
    .A2(_05088_),
    .B1(net954),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00006_));
 sky130_fd_sc_hd__nand2_1 _09057_ (.A(_03391_),
    .B(_04255_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05089_));
 sky130_fd_sc_hd__nor2_1 _09058_ (.A(_02859_),
    .B(_04257_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05090_));
 sky130_fd_sc_hd__or2_1 _09059_ (.A(_02859_),
    .B(_04257_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05091_));
 sky130_fd_sc_hd__a22o_1 _09060_ (.A1(net1588),
    .A2(_05089_),
    .B1(_05090_),
    .B2(net1542),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00026_));
 sky130_fd_sc_hd__o31a_1 _09061_ (.A1(net424),
    .A2(_02969_),
    .A3(_02995_),
    .B1(net523),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05092_));
 sky130_fd_sc_hd__a31o_1 _09062_ (.A1(net463),
    .A2(_04191_),
    .A3(_04556_),
    .B1(_05092_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00005_));
 sky130_fd_sc_hd__nor2_1 _09063_ (.A(net447),
    .B(net455),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05093_));
 sky130_fd_sc_hd__or2_1 _09064_ (.A(net447),
    .B(net458),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05094_));
 sky130_fd_sc_hd__a211o_1 _09065_ (.A1(net444),
    .A2(net455),
    .B1(_03013_),
    .C1(_05093_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05095_));
 sky130_fd_sc_hd__a32o_1 _09066_ (.A1(net439),
    .A2(\top.sram_interface.word_cnt[9] ),
    .A3(_05094_),
    .B1(_05095_),
    .B2(net1581),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00049_));
 sky130_fd_sc_hd__nor2_2 _09067_ (.A(_03013_),
    .B(_05094_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05096_));
 sky130_fd_sc_hd__a21o_1 _09068_ (.A1(net443),
    .A2(net450),
    .B1(_05096_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05097_));
 sky130_fd_sc_hd__nand2_1 _09069_ (.A(net460),
    .B(net526),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05098_));
 sky130_fd_sc_hd__a32o_1 _09070_ (.A1(net462),
    .A2(net526),
    .A3(_02910_),
    .B1(_05097_),
    .B2(net546),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05099_));
 sky130_fd_sc_hd__or3b_1 _09071_ (.A(_02715_),
    .B(_05099_),
    .C_N(_02915_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00038_));
 sky130_fd_sc_hd__or3_1 _09072_ (.A(net447),
    .B(_02562_),
    .C(_03013_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05100_));
 sky130_fd_sc_hd__a22o_1 _09073_ (.A1(net457),
    .A2(net1040),
    .B1(_05100_),
    .B2(net1237),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00050_));
 sky130_fd_sc_hd__nor2_1 _09074_ (.A(_02796_),
    .B(_02799_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05101_));
 sky130_fd_sc_hd__a32o_1 _09075_ (.A1(net452),
    .A2(_02916_),
    .A3(_02922_),
    .B1(_02900_),
    .B2(net466),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05102_));
 sky130_fd_sc_hd__o31a_1 _09076_ (.A1(_02794_),
    .A2(_05101_),
    .A3(_05102_),
    .B1(net542),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05103_));
 sky130_fd_sc_hd__a221o_1 _09077_ (.A1(net458),
    .A2(net545),
    .B1(\top.sram_interface.word_cnt[2] ),
    .B2(net446),
    .C1(_02590_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05104_));
 sky130_fd_sc_hd__a31o_1 _09078_ (.A1(net455),
    .A2(\top.sram_interface.word_cnt[7] ),
    .A3(_02797_),
    .B1(_05104_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05105_));
 sky130_fd_sc_hd__a21o_1 _09079_ (.A1(net442),
    .A2(net451),
    .B1(_05096_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05106_));
 sky130_fd_sc_hd__a211o_1 _09080_ (.A1(net533),
    .A2(_05106_),
    .B1(_05105_),
    .C1(_05103_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00051_));
 sky130_fd_sc_hd__a21o_1 _09081_ (.A1(net443),
    .A2(net459),
    .B1(_05096_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05107_));
 sky130_fd_sc_hd__a21o_1 _09082_ (.A1(net443),
    .A2(net450),
    .B1(_05107_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05108_));
 sky130_fd_sc_hd__o21a_1 _09083_ (.A1(net451),
    .A2(_05108_),
    .B1(\top.sram_interface.word_cnt[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05109_));
 sky130_fd_sc_hd__a221o_1 _09084_ (.A1(net460),
    .A2(\top.sram_interface.word_cnt[2] ),
    .B1(net356),
    .B2(\top.hTree.write_HT_fin ),
    .C1(_05109_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05110_));
 sky130_fd_sc_hd__a31o_1 _09085_ (.A1(net459),
    .A2(net534),
    .A3(_02576_),
    .B1(_05110_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00052_));
 sky130_fd_sc_hd__a221o_1 _09086_ (.A1(\top.sram_interface.word_cnt[6] ),
    .A2(_02795_),
    .B1(_02839_),
    .B2(net537),
    .C1(_05076_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05111_));
 sky130_fd_sc_hd__and4b_1 _09087_ (.A_N(\top.sram_interface.CB_write_counter[1] ),
    .B(\top.sram_interface.CB_write_counter[0] ),
    .C(net460),
    .D(\top.sram_interface.word_cnt[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05112_));
 sky130_fd_sc_hd__a211o_1 _09088_ (.A1(net527),
    .A2(_05107_),
    .B1(_05111_),
    .C1(_05112_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00039_));
 sky130_fd_sc_hd__a22o_1 _09089_ (.A1(net455),
    .A2(\top.sram_interface.word_cnt[4] ),
    .B1(_05100_),
    .B2(net1040),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00040_));
 sky130_fd_sc_hd__a31o_1 _09090_ (.A1(\top.sram_interface.CB_write_counter[1] ),
    .A2(\top.sram_interface.CB_write_counter[0] ),
    .A3(net460),
    .B1(_05107_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05113_));
 sky130_fd_sc_hd__or4b_1 _09091_ (.A(\top.sram_interface.TRN_counter[2] ),
    .B(\top.sram_interface.TRN_counter[1] ),
    .C(\top.sram_interface.TRN_counter[0] ),
    .D_N(net452),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05114_));
 sky130_fd_sc_hd__o21ai_1 _09092_ (.A1(net442),
    .A2(net423),
    .B1(_05114_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05115_));
 sky130_fd_sc_hd__a22o_1 _09093_ (.A1(net526),
    .A2(_05113_),
    .B1(_05115_),
    .B2(net536),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05116_));
 sky130_fd_sc_hd__a221o_1 _09094_ (.A1(net456),
    .A2(\top.sram_interface.word_cnt[2] ),
    .B1(net527),
    .B2(net447),
    .C1(_05116_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00041_));
 sky130_fd_sc_hd__o21a_1 _09095_ (.A1(_03013_),
    .A2(_05093_),
    .B1(\top.sram_interface.word_cnt[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05117_));
 sky130_fd_sc_hd__a221o_1 _09096_ (.A1(net447),
    .A2(net1581),
    .B1(net527),
    .B2(_02795_),
    .C1(_05117_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00042_));
 sky130_fd_sc_hd__a211o_1 _09097_ (.A1(net443),
    .A2(net462),
    .B1(net451),
    .C1(_05107_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05118_));
 sky130_fd_sc_hd__a22o_1 _09098_ (.A1(net546),
    .A2(_02839_),
    .B1(_05118_),
    .B2(\top.sram_interface.word_cnt[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05119_));
 sky130_fd_sc_hd__a32o_1 _09099_ (.A1(net462),
    .A2(net534),
    .A3(_02582_),
    .B1(_03038_),
    .B2(_02575_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05120_));
 sky130_fd_sc_hd__or2_1 _09100_ (.A(_05119_),
    .B(_05120_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00043_));
 sky130_fd_sc_hd__nand2_1 _09101_ (.A(\top.hTree.wait_cnt ),
    .B(net255),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05121_));
 sky130_fd_sc_hd__a32o_1 _09102_ (.A1(\top.hTree.wait_cnt ),
    .A2(net1522),
    .A3(net254),
    .B1(_05091_),
    .B2(net1542),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00027_));
 sky130_fd_sc_hd__mux2_1 _09103_ (.A0(net1004),
    .A1(net1604),
    .S(net254),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00018_));
 sky130_fd_sc_hd__or2_2 _09104_ (.A(\top.histogram.init_edge ),
    .B(_05080_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05122_));
 sky130_fd_sc_hd__nor2_1 _09105_ (.A(net481),
    .B(_05122_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05123_));
 sky130_fd_sc_hd__nor2_1 _09106_ (.A(_02594_),
    .B(_05122_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05124_));
 sky130_fd_sc_hd__or2_1 _09107_ (.A(_02594_),
    .B(_05122_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05125_));
 sky130_fd_sc_hd__nand2_1 _09108_ (.A(net453),
    .B(_05125_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05126_));
 sky130_fd_sc_hd__and4b_1 _09109_ (.A_N(\top.histogram.out_of_init ),
    .B(\top.histogram.eof_n ),
    .C(_02561_),
    .D(_05124_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05127_));
 sky130_fd_sc_hd__and3_1 _09110_ (.A(net439),
    .B(\top.histogram.state[7] ),
    .C(_05124_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05128_));
 sky130_fd_sc_hd__a211o_1 _09111_ (.A1(\top.histogram.state[0] ),
    .A2(_05126_),
    .B1(_05127_),
    .C1(_05128_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00028_));
 sky130_fd_sc_hd__nor2_1 _09112_ (.A(_03369_),
    .B(_05122_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05129_));
 sky130_fd_sc_hd__a22o_1 _09113_ (.A1(_02417_),
    .A2(net1750),
    .B1(_05129_),
    .B2(_02416_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00029_));
 sky130_fd_sc_hd__a21o_1 _09114_ (.A1(net444),
    .A2(_05124_),
    .B1(_02417_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05130_));
 sky130_fd_sc_hd__a22o_1 _09115_ (.A1(_05079_),
    .A2(_05124_),
    .B1(_05130_),
    .B2(net1446),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00030_));
 sky130_fd_sc_hd__a22o_1 _09116_ (.A1(net353),
    .A2(_05123_),
    .B1(_05130_),
    .B2(net1658),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00031_));
 sky130_fd_sc_hd__and4b_1 _09117_ (.A_N(_03368_),
    .B(_05124_),
    .C(\top.histogram.eof_n ),
    .D(\top.dut.out_valid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05131_));
 sky130_fd_sc_hd__a221o_1 _09118_ (.A1(_02417_),
    .A2(\top.histogram.eof_n ),
    .B1(net360),
    .B2(_05122_),
    .C1(_05131_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00032_));
 sky130_fd_sc_hd__a21o_1 _09119_ (.A1(net453),
    .A2(\top.histogram.state[1] ),
    .B1(net1786),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05132_));
 sky130_fd_sc_hd__and2_1 _09120_ (.A(_05126_),
    .B(_05132_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00033_));
 sky130_fd_sc_hd__a211o_1 _09121_ (.A1(\top.histogram.init_edge ),
    .A2(_02416_),
    .B1(_03244_),
    .C1(_05080_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05133_));
 sky130_fd_sc_hd__nand2_1 _09122_ (.A(_02610_),
    .B(_05133_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05134_));
 sky130_fd_sc_hd__a21o_1 _09123_ (.A1(_02417_),
    .A2(net1514),
    .B1(_05134_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00034_));
 sky130_fd_sc_hd__a22o_1 _09124_ (.A1(\top.histogram.state[6] ),
    .A2(_05124_),
    .B1(_05130_),
    .B2(net1479),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00035_));
 sky130_fd_sc_hd__or4_1 _09125_ (.A(\top.histogram.state[7] ),
    .B(\top.histogram.state[3] ),
    .C(\top.histogram.state[5] ),
    .D(\top.histogram.state[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05135_));
 sky130_fd_sc_hd__or4_1 _09126_ (.A(\top.histogram.eof_n ),
    .B(\top.histogram.state[0] ),
    .C(\top.histogram.state[2] ),
    .D(\top.histogram.state[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05136_));
 sky130_fd_sc_hd__or3_1 _09127_ (.A(_05125_),
    .B(_05135_),
    .C(_05136_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05137_));
 sky130_fd_sc_hd__or4b_1 _09128_ (.A(_02417_),
    .B(_05127_),
    .C(_05131_),
    .D_N(_05137_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05138_));
 sky130_fd_sc_hd__a22o_1 _09129_ (.A1(net360),
    .A2(_05122_),
    .B1(_05138_),
    .B2(net1574),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00036_));
 sky130_fd_sc_hd__a21o_1 _09130_ (.A1(net1517),
    .A2(_05138_),
    .B1(_05134_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00037_));
 sky130_fd_sc_hd__o211a_1 _09131_ (.A1(\top.sram_interface.word_cnt[9] ),
    .A2(net545),
    .B1(_02587_),
    .C1(net460),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05139_));
 sky130_fd_sc_hd__and2b_1 _09132_ (.A_N(_02906_),
    .B(_02795_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05140_));
 sky130_fd_sc_hd__a32o_1 _09133_ (.A1(net455),
    .A2(\top.sram_interface.word_cnt[7] ),
    .A3(_02798_),
    .B1(_05096_),
    .B2(net542),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05141_));
 sky130_fd_sc_hd__or3_1 _09134_ (.A(_05139_),
    .B(_05140_),
    .C(_05141_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05142_));
 sky130_fd_sc_hd__or4b_1 _09135_ (.A(_02862_),
    .B(_05142_),
    .C(net304),
    .D_N(_02585_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05143_));
 sky130_fd_sc_hd__and4bb_1 _09136_ (.A_N(\top.findLeastValue.histo_index[8] ),
    .B_N(_02575_),
    .C(_02816_),
    .D(\top.sram_interface.zero_cnt[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05144_));
 sky130_fd_sc_hd__a31o_1 _09137_ (.A1(net443),
    .A2(_02817_),
    .A3(_05144_),
    .B1(_03391_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05145_));
 sky130_fd_sc_hd__or4_1 _09138_ (.A(_02858_),
    .B(_02880_),
    .C(_05143_),
    .D(_05145_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05146_));
 sky130_fd_sc_hd__a41o_1 _09139_ (.A1(net543),
    .A2(net452),
    .A3(_02916_),
    .A4(_02921_),
    .B1(_05146_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05147_));
 sky130_fd_sc_hd__a311o_1 _09140_ (.A1(net543),
    .A2(net466),
    .A3(_02901_),
    .B1(_05147_),
    .C1(_02802_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00044_));
 sky130_fd_sc_hd__o211a_1 _09141_ (.A1(\top.WorR ),
    .A2(_02856_),
    .B1(_02852_),
    .C1(net448),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05148_));
 sky130_fd_sc_hd__a2bb2o_1 _09142_ (.A1_N(_02840_),
    .A2_N(_03390_),
    .B1(_05148_),
    .B2(_02845_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05149_));
 sky130_fd_sc_hd__o211a_1 _09143_ (.A1(net462),
    .A2(net456),
    .B1(\top.sram_interface.word_cnt[14] ),
    .C1(net439),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05150_));
 sky130_fd_sc_hd__o21a_1 _09144_ (.A1(net451),
    .A2(_05096_),
    .B1(\top.sram_interface.word_cnt[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05151_));
 sky130_fd_sc_hd__a221o_1 _09145_ (.A1(net448),
    .A2(_02860_),
    .B1(_05149_),
    .B2(net544),
    .C1(_05151_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05152_));
 sky130_fd_sc_hd__or2_1 _09146_ (.A(_05150_),
    .B(_05152_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00045_));
 sky130_fd_sc_hd__a21oi_1 _09147_ (.A1(net457),
    .A2(net361),
    .B1(_02596_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05153_));
 sky130_fd_sc_hd__o311a_1 _09148_ (.A1(\top.sram_interface.CB_write_counter[1] ),
    .A2(\top.sram_interface.CB_write_counter[0] ),
    .A3(_05098_),
    .B1(_05153_),
    .C1(net317),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05154_));
 sky130_fd_sc_hd__a21bo_1 _09149_ (.A1(net537),
    .A2(_05108_),
    .B1_N(_05154_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00046_));
 sky130_fd_sc_hd__a22o_1 _09150_ (.A1(net455),
    .A2(\top.sram_interface.word_cnt[13] ),
    .B1(_05100_),
    .B2(net1047),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00047_));
 sky130_fd_sc_hd__and3b_1 _09151_ (.A_N(_05144_),
    .B(net456),
    .C(net443),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05155_));
 sky130_fd_sc_hd__a221o_1 _09152_ (.A1(net442),
    .A2(net462),
    .B1(net451),
    .B2(\top.sram_interface.TRN_counter[2] ),
    .C1(_05096_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05156_));
 sky130_fd_sc_hd__o21a_1 _09153_ (.A1(_05155_),
    .A2(_05156_),
    .B1(net536),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05157_));
 sky130_fd_sc_hd__a22o_1 _09154_ (.A1(net440),
    .A2(net451),
    .B1(net456),
    .B2(net406),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05158_));
 sky130_fd_sc_hd__a221o_1 _09155_ (.A1(net447),
    .A2(\top.sram_interface.word_cnt[14] ),
    .B1(_05158_),
    .B2(net535),
    .C1(_02607_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05159_));
 sky130_fd_sc_hd__or2_1 _09156_ (.A(_05157_),
    .B(_05159_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00048_));
 sky130_fd_sc_hd__a31o_1 _09157_ (.A1(\top.cb_syn.curr_state[0] ),
    .A2(_04206_),
    .A3(_04546_),
    .B1(_04544_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00003_));
 sky130_fd_sc_hd__and4b_1 _09158_ (.A_N(\top.cb_syn.char_path_n[2] ),
    .B(net516),
    .C(net463),
    .D(_04562_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05160_));
 sky130_fd_sc_hd__o31a_1 _09159_ (.A1(\top.cb_syn.pulse_first ),
    .A2(net424),
    .A3(_02890_),
    .B1(net522),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05161_));
 sky130_fd_sc_hd__or3_1 _09160_ (.A(_04557_),
    .B(_05160_),
    .C(_05161_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00007_));
 sky130_fd_sc_hd__o21a_1 _09161_ (.A1(\top.cb_syn.end_check ),
    .A2(net424),
    .B1(\top.cb_syn.curr_state[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05162_));
 sky130_fd_sc_hd__a22oi_1 _09162_ (.A1(net525),
    .A2(_04551_),
    .B1(_04606_),
    .B2(net520),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05163_));
 sky130_fd_sc_hd__nor2_1 _09163_ (.A(_04206_),
    .B(_05163_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05164_));
 sky130_fd_sc_hd__or3_1 _09164_ (.A(_04547_),
    .B(_05162_),
    .C(_05164_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00008_));
 sky130_fd_sc_hd__or3b_1 _09165_ (.A(net424),
    .B(_02890_),
    .C_N(_05084_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05165_));
 sky130_fd_sc_hd__and4b_1 _09166_ (.A_N(\top.cb_syn.char_path_n[1] ),
    .B(net515),
    .C(net464),
    .D(_04201_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05166_));
 sky130_fd_sc_hd__and4b_1 _09167_ (.A_N(_02969_),
    .B(_02993_),
    .C(\top.cb_syn.curr_state[2] ),
    .D(net464),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05167_));
 sky130_fd_sc_hd__a211o_1 _09168_ (.A1(net519),
    .A2(_05165_),
    .B1(_05166_),
    .C1(_05167_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00009_));
 sky130_fd_sc_hd__or3b_1 _09169_ (.A(\top.cb_syn.setup ),
    .B(net488),
    .C_N(\top.cb_syn.curr_state[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05168_));
 sky130_fd_sc_hd__a21bo_1 _09170_ (.A1(net488),
    .A2(net524),
    .B1_N(_05168_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05169_));
 sky130_fd_sc_hd__a22o_1 _09171_ (.A1(_02581_),
    .A2(_02887_),
    .B1(_04605_),
    .B2(_02551_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05170_));
 sky130_fd_sc_hd__o31a_1 _09172_ (.A1(_02896_),
    .A2(_05169_),
    .A3(_05170_),
    .B1(net464),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05171_));
 sky130_fd_sc_hd__a221o_1 _09173_ (.A1(net524),
    .A2(net424),
    .B1(_04585_),
    .B2(_05086_),
    .C1(_05171_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00004_));
 sky130_fd_sc_hd__a22o_1 _09174_ (.A1(net1378),
    .A2(_02567_),
    .B1(\top.WB.curr_state[0] ),
    .B2(_02615_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00002_));
 sky130_fd_sc_hd__a22o_1 _09175_ (.A1(\top.WB.curr_state[1] ),
    .A2(_02567_),
    .B1(\top.WB.curr_state[0] ),
    .B2(_02617_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00001_));
 sky130_fd_sc_hd__o21ai_1 _09176_ (.A1(_02567_),
    .A2(_02572_),
    .B1(_02618_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_00000_));
 sky130_fd_sc_hd__a22o_1 _09177_ (.A1(net1511),
    .A2(_05054_),
    .B1(_05090_),
    .B2(\top.hTree.state[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00025_));
 sky130_fd_sc_hd__nor4_1 _09178_ (.A(\top.controller.fin_reg[1] ),
    .B(\top.controller.fin_reg[2] ),
    .C(\top.controller.fin_reg[3] ),
    .D(\top.controller.fin_reg[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05172_));
 sky130_fd_sc_hd__and3_1 _09179_ (.A(net1592),
    .B(\top.controller.fin_reg[7] ),
    .C(_05172_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00013_));
 sky130_fd_sc_hd__a32o_1 _09180_ (.A1(net1699),
    .A2(\top.hTree.state[2] ),
    .A3(net254),
    .B1(_05091_),
    .B2(\top.hTree.state[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00024_));
 sky130_fd_sc_hd__o21a_1 _09181_ (.A1(_02514_),
    .A2(_02835_),
    .B1(\top.hTree.write_HT_fin ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05173_));
 sky130_fd_sc_hd__and3_1 _09182_ (.A(net287),
    .B(_05050_),
    .C(_05173_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05174_));
 sky130_fd_sc_hd__or3_1 _09183_ (.A(net248),
    .B(_05058_),
    .C(_05174_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05175_));
 sky130_fd_sc_hd__a22o_1 _09184_ (.A1(net1004),
    .A2(net254),
    .B1(_05175_),
    .B2(net470),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00017_));
 sky130_fd_sc_hd__a22o_1 _09185_ (.A1(\top.hTree.state[4] ),
    .A2(net255),
    .B1(_05121_),
    .B2(net1522),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00023_));
 sky130_fd_sc_hd__mux2_1 _09186_ (.A0(net1677),
    .A1(_05051_),
    .S(net254),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00022_));
 sky130_fd_sc_hd__mux2_1 _09187_ (.A0(\top.hTree.state[3] ),
    .A1(_05057_),
    .S(net256),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05176_));
 sky130_fd_sc_hd__or2_1 _09188_ (.A(_02866_),
    .B(_05176_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00021_));
 sky130_fd_sc_hd__a22o_1 _09189_ (.A1(\top.hTree.state[3] ),
    .A2(net254),
    .B1(_05121_),
    .B2(net1637),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00020_));
 sky130_fd_sc_hd__a22o_1 _09190_ (.A1(_02851_),
    .A2(_04255_),
    .B1(_05173_),
    .B2(net470),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05177_));
 sky130_fd_sc_hd__a22o_1 _09191_ (.A1(net1604),
    .A2(_04257_),
    .B1(_05177_),
    .B2(_03393_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00019_));
 sky130_fd_sc_hd__mux2_1 _09192_ (.A0(net514),
    .A1(_02888_),
    .S(net463),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05178_));
 sky130_fd_sc_hd__a21o_1 _09193_ (.A1(_04542_),
    .A2(_04543_),
    .B1(_05178_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00011_));
 sky130_fd_sc_hd__o211a_1 _09194_ (.A1(\top.cb_syn.char_path_n[1] ),
    .A2(_04201_),
    .B1(_04563_),
    .C1(net463),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05179_));
 sky130_fd_sc_hd__o22ai_1 _09195_ (.A1(_04541_),
    .A2(_04548_),
    .B1(_05179_),
    .B2(_02543_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_00010_));
 sky130_fd_sc_hd__or4bb_1 _09196_ (.A(\top.controller.fin_reg[1] ),
    .B(\top.controller.fin_reg[4] ),
    .C_N(\top.controller.fin_reg[3] ),
    .D_N(\top.controller.fin_reg[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05180_));
 sky130_fd_sc_hd__nand3_1 _09197_ (.A(\top.controller.fin_reg[5] ),
    .B(\top.controller.fin_reg[6] ),
    .C(\top.controller.fin_reg[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05181_));
 sky130_fd_sc_hd__nor2_1 _09198_ (.A(_05180_),
    .B(_05181_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_00015_));
 sky130_fd_sc_hd__or4b_1 _09199_ (.A(net1778),
    .B(\top.controller.fin_reg[2] ),
    .C(\top.controller.fin_reg[4] ),
    .D_N(\top.controller.fin_reg[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05182_));
 sky130_fd_sc_hd__nor2_1 _09200_ (.A(_05181_),
    .B(_05182_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_00012_));
 sky130_fd_sc_hd__or4_1 _09201_ (.A(\top.controller.fin_reg[1] ),
    .B(\top.controller.fin_reg[2] ),
    .C(net1681),
    .D(\top.controller.fin_reg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05183_));
 sky130_fd_sc_hd__nor2_1 _09202_ (.A(_05181_),
    .B(_05183_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_00016_));
 sky130_fd_sc_hd__or4b_1 _09203_ (.A(net1679),
    .B(_05183_),
    .C(net1592),
    .D_N(\top.controller.fin_reg[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05184_));
 sky130_fd_sc_hd__inv_2 _09204_ (.A(_05184_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_00014_));
 sky130_fd_sc_hd__nor3b_1 _09205_ (.A(\top.header_synthesis.start ),
    .B(_03375_),
    .C_N(_03372_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05185_));
 sky130_fd_sc_hd__inv_2 _09206_ (.A(_05185_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05186_));
 sky130_fd_sc_hd__or4_1 _09207_ (.A(\top.cb_syn.num_lefts[5] ),
    .B(\top.cb_syn.num_lefts[4] ),
    .C(\top.cb_syn.num_lefts[3] ),
    .D(\top.cb_syn.num_lefts[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05187_));
 sky130_fd_sc_hd__o41a_1 _09208_ (.A1(\top.cb_syn.num_lefts[7] ),
    .A2(\top.cb_syn.num_lefts[6] ),
    .A3(_04604_),
    .A4(_05187_),
    .B1(_02566_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05188_));
 sky130_fd_sc_hd__a32o_1 _09209_ (.A1(net1085),
    .A2(net291),
    .A3(_05188_),
    .B1(\top.header_synthesis.write_num_lefts ),
    .B2(_03375_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\top.header_synthesis.next_write_num_lefts ));
 sky130_fd_sc_hd__o221a_1 _09210_ (.A1(net491),
    .A2(\top.header_synthesis.write_char_path ),
    .B1(_03382_),
    .B2(_02566_),
    .C1(_05186_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\top.header_synthesis.next_write_char_path ));
 sky130_fd_sc_hd__a21o_1 _09211_ (.A1(_02956_),
    .A2(_02964_),
    .B1(_02961_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05189_));
 sky130_fd_sc_hd__o221a_1 _09212_ (.A1(_02529_),
    .A2(\top.cb_syn.zero_count[4] ),
    .B1(_02958_),
    .B2(_02959_),
    .C1(_05189_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05190_));
 sky130_fd_sc_hd__o21bai_1 _09213_ (.A1(_02954_),
    .A2(_05190_),
    .B1_N(_02957_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05191_));
 sky130_fd_sc_hd__a21oi_1 _09214_ (.A1(_02955_),
    .A2(_05191_),
    .B1(_02962_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05192_));
 sky130_fd_sc_hd__or3_1 _09215_ (.A(_02963_),
    .B(_02968_),
    .C(_05192_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05193_));
 sky130_fd_sc_hd__inv_2 _09216_ (.A(_05193_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05194_));
 sky130_fd_sc_hd__a211o_1 _09217_ (.A1(\top.header_synthesis.write_zeroes ),
    .A2(_05193_),
    .B1(net491),
    .C1(_02565_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05195_));
 sky130_fd_sc_hd__a311o_1 _09218_ (.A1(_03371_),
    .A2(_03388_),
    .A3(_05195_),
    .B1(net291),
    .C1(\top.header_synthesis.write_num_lefts ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05196_));
 sky130_fd_sc_hd__a21bo_1 _09219_ (.A1(\top.header_synthesis.write_num_lefts ),
    .A2(_03375_),
    .B1_N(_05196_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\top.header_synthesis.next_enable ));
 sky130_fd_sc_hd__o21a_1 _09220_ (.A1(net491),
    .A2(net1704),
    .B1(_03371_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\top.header_synthesis.next_start ));
 sky130_fd_sc_hd__nor2_1 _09221_ (.A(net490),
    .B(net1674),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05197_));
 sky130_fd_sc_hd__o21ai_1 _09222_ (.A1(_03372_),
    .A2(_05197_),
    .B1(_03376_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\top.header_synthesis.next_char_added ));
 sky130_fd_sc_hd__mux2_1 _09223_ (.A0(\top.header_synthesis.header[0] ),
    .A1(\top.cb_syn.char_index[0] ),
    .S(net490),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05198_));
 sky130_fd_sc_hd__and2_1 _09224_ (.A(net296),
    .B(_05198_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\top.header_synthesis.next_header[0] ));
 sky130_fd_sc_hd__mux2_1 _09225_ (.A0(\top.header_synthesis.header[1] ),
    .A1(\top.cb_syn.char_index[1] ),
    .S(net490),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05199_));
 sky130_fd_sc_hd__mux2_1 _09226_ (.A0(net1408),
    .A1(_05199_),
    .S(net296),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\top.header_synthesis.next_header[1] ));
 sky130_fd_sc_hd__mux2_1 _09227_ (.A0(\top.header_synthesis.header[2] ),
    .A1(\top.cb_syn.char_index[2] ),
    .S(net490),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05200_));
 sky130_fd_sc_hd__mux2_1 _09228_ (.A0(net1081),
    .A1(_05200_),
    .S(net296),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\top.header_synthesis.next_header[2] ));
 sky130_fd_sc_hd__mux2_1 _09229_ (.A0(\top.header_synthesis.header[3] ),
    .A1(\top.cb_syn.char_index[3] ),
    .S(net490),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05201_));
 sky130_fd_sc_hd__mux2_1 _09230_ (.A0(net1147),
    .A1(_05201_),
    .S(net296),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\top.header_synthesis.next_header[3] ));
 sky130_fd_sc_hd__mux2_1 _09231_ (.A0(\top.header_synthesis.header[4] ),
    .A1(\top.cb_syn.char_index[4] ),
    .S(net490),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05202_));
 sky130_fd_sc_hd__mux2_1 _09232_ (.A0(net1173),
    .A1(_05202_),
    .S(net296),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\top.header_synthesis.next_header[4] ));
 sky130_fd_sc_hd__mux2_1 _09233_ (.A0(\top.header_synthesis.header[5] ),
    .A1(\top.cb_syn.char_index[5] ),
    .S(net490),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05203_));
 sky130_fd_sc_hd__mux2_1 _09234_ (.A0(net1083),
    .A1(_05203_),
    .S(net296),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\top.header_synthesis.next_header[5] ));
 sky130_fd_sc_hd__mux2_1 _09235_ (.A0(\top.header_synthesis.header[6] ),
    .A1(\top.cb_syn.char_index[6] ),
    .S(net490),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05204_));
 sky130_fd_sc_hd__mux2_1 _09236_ (.A0(net1247),
    .A1(_05204_),
    .S(net296),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\top.header_synthesis.next_header[6] ));
 sky130_fd_sc_hd__mux2_1 _09237_ (.A0(\top.header_synthesis.header[7] ),
    .A1(\top.cb_syn.char_index[7] ),
    .S(net490),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05205_));
 sky130_fd_sc_hd__mux2_1 _09238_ (.A0(net1064),
    .A1(_05205_),
    .S(net296),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\top.header_synthesis.next_header[7] ));
 sky130_fd_sc_hd__or2_1 _09239_ (.A(net490),
    .B(\top.header_synthesis.header[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05206_));
 sky130_fd_sc_hd__mux2_1 _09240_ (.A0(net1232),
    .A1(_05206_),
    .S(net296),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\top.header_synthesis.next_header[8] ));
 sky130_fd_sc_hd__and3_2 _09241_ (.A(\top.header_synthesis.write_zeroes ),
    .B(_03388_),
    .C(_05194_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05207_));
 sky130_fd_sc_hd__a21oi_4 _09242_ (.A1(\top.header_synthesis.write_zeroes ),
    .A2(_03388_),
    .B1(net491),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05208_));
 sky130_fd_sc_hd__mux2_1 _09243_ (.A0(_05207_),
    .A1(_05208_),
    .S(\top.cb_syn.zero_count[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\top.header_synthesis.next_zero_count[0] ));
 sky130_fd_sc_hd__nand2_1 _09244_ (.A(\top.cb_syn.zero_count[0] ),
    .B(\top.cb_syn.zero_count[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05209_));
 sky130_fd_sc_hd__or2_1 _09245_ (.A(\top.cb_syn.zero_count[0] ),
    .B(\top.cb_syn.zero_count[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05210_));
 sky130_fd_sc_hd__a32o_1 _09246_ (.A1(_05207_),
    .A2(_05209_),
    .A3(_05210_),
    .B1(_05208_),
    .B2(net1713),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\top.header_synthesis.next_zero_count[1] ));
 sky130_fd_sc_hd__nand2_1 _09247_ (.A(_02558_),
    .B(_05209_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05211_));
 sky130_fd_sc_hd__or2_1 _09248_ (.A(_02558_),
    .B(_05209_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05212_));
 sky130_fd_sc_hd__a32o_1 _09249_ (.A1(_05207_),
    .A2(_05211_),
    .A3(_05212_),
    .B1(_05208_),
    .B2(net1605),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\top.header_synthesis.next_zero_count[2] ));
 sky130_fd_sc_hd__nand2_1 _09250_ (.A(_02557_),
    .B(_05212_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05213_));
 sky130_fd_sc_hd__nor2_1 _09251_ (.A(_02557_),
    .B(_05212_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05214_));
 sky130_fd_sc_hd__inv_2 _09252_ (.A(_05214_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05215_));
 sky130_fd_sc_hd__a32o_1 _09253_ (.A1(_05207_),
    .A2(_05213_),
    .A3(_05215_),
    .B1(_05208_),
    .B2(net1561),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\top.header_synthesis.next_zero_count[3] ));
 sky130_fd_sc_hd__nand2_1 _09254_ (.A(\top.cb_syn.zero_count[4] ),
    .B(_05214_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05216_));
 sky130_fd_sc_hd__or2_1 _09255_ (.A(\top.cb_syn.zero_count[4] ),
    .B(_05214_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05217_));
 sky130_fd_sc_hd__a32o_1 _09256_ (.A1(_05207_),
    .A2(_05216_),
    .A3(_05217_),
    .B1(_05208_),
    .B2(\top.cb_syn.zero_count[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\top.header_synthesis.next_zero_count[4] ));
 sky130_fd_sc_hd__nor2_1 _09257_ (.A(_02559_),
    .B(_05216_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05218_));
 sky130_fd_sc_hd__inv_2 _09258_ (.A(_05218_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05219_));
 sky130_fd_sc_hd__nand2_1 _09259_ (.A(_02559_),
    .B(_05216_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05220_));
 sky130_fd_sc_hd__a32o_1 _09260_ (.A1(_05207_),
    .A2(_05219_),
    .A3(_05220_),
    .B1(_05208_),
    .B2(net1642),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\top.header_synthesis.next_zero_count[5] ));
 sky130_fd_sc_hd__or2_1 _09261_ (.A(\top.cb_syn.zero_count[6] ),
    .B(_05218_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05221_));
 sky130_fd_sc_hd__nand2_1 _09262_ (.A(\top.cb_syn.zero_count[6] ),
    .B(_05218_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05222_));
 sky130_fd_sc_hd__a32o_1 _09263_ (.A1(_05207_),
    .A2(_05221_),
    .A3(_05222_),
    .B1(_05208_),
    .B2(net1708),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\top.header_synthesis.next_zero_count[6] ));
 sky130_fd_sc_hd__a21o_1 _09264_ (.A1(_05207_),
    .A2(_05222_),
    .B1(_05208_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05223_));
 sky130_fd_sc_hd__nor2_1 _09265_ (.A(\top.cb_syn.zero_count[7] ),
    .B(_05222_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05224_));
 sky130_fd_sc_hd__a22o_1 _09266_ (.A1(net1666),
    .A2(_05223_),
    .B1(_05224_),
    .B2(_05207_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\top.header_synthesis.next_zero_count[7] ));
 sky130_fd_sc_hd__o31a_1 _09267_ (.A1(net1684),
    .A2(_04046_),
    .A3(\top.dut.bits_in_buf_next[0] ),
    .B1(_04098_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\top.dut.bit_buf_next[0] ));
 sky130_fd_sc_hd__o21a_1 _09268_ (.A1(_04046_),
    .A2(\top.dut.bits_in_buf_next[1] ),
    .B1(_04094_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\top.dut.bit_buf_next[1] ));
 sky130_fd_sc_hd__o21a_1 _09269_ (.A1(_04046_),
    .A2(_04067_),
    .B1(_04090_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\top.dut.bit_buf_next[2] ));
 sky130_fd_sc_hd__and2_1 _09270_ (.A(_04046_),
    .B(_04086_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\top.dut.bit_buf_next[3] ));
 sky130_fd_sc_hd__nor2_1 _09271_ (.A(_04044_),
    .B(_04095_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05225_));
 sky130_fd_sc_hd__o21a_1 _09272_ (.A1(net343),
    .A2(_05225_),
    .B1(_04081_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\top.dut.bit_buf_next[4] ));
 sky130_fd_sc_hd__o21a_1 _09273_ (.A1(net343),
    .A2(_04067_),
    .B1(_04046_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05226_));
 sky130_fd_sc_hd__o21a_1 _09274_ (.A1(_04057_),
    .A2(_05226_),
    .B1(_04076_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\top.dut.bit_buf_next[5] ));
 sky130_fd_sc_hd__and2_1 _09275_ (.A(_04072_),
    .B(_05226_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\top.dut.bit_buf_next[6] ));
 sky130_fd_sc_hd__and2_1 _09276_ (.A(net343),
    .B(_04054_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\top.dut.bit_buf_next[7] ));
 sky130_fd_sc_hd__and2_1 _09277_ (.A(net344),
    .B(_04053_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\top.dut.bit_buf_next[8] ));
 sky130_fd_sc_hd__and2_1 _09278_ (.A(net343),
    .B(_04051_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\top.dut.bit_buf_next[9] ));
 sky130_fd_sc_hd__and2_1 _09279_ (.A(net344),
    .B(_04050_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\top.dut.bit_buf_next[10] ));
 sky130_fd_sc_hd__and2_1 _09280_ (.A(net343),
    .B(_04063_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\top.dut.bit_buf_next[11] ));
 sky130_fd_sc_hd__and2_1 _09281_ (.A(net343),
    .B(_04062_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\top.dut.bit_buf_next[12] ));
 sky130_fd_sc_hd__and2_1 _09282_ (.A(net343),
    .B(_04058_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\top.dut.bit_buf_next[13] ));
 sky130_fd_sc_hd__and4b_1 _09283_ (.A_N(\top.translation.totalEn ),
    .B(_05023_),
    .C(_05024_),
    .D(\top.translation.writeEn ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05227_));
 sky130_fd_sc_hd__mux4_1 _09284_ (.A0(\top.histogram.total[20] ),
    .A1(\top.histogram.total[21] ),
    .A2(\top.histogram.total[22] ),
    .A3(\top.histogram.total[23] ),
    .S0(net508),
    .S1(net506),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05228_));
 sky130_fd_sc_hd__mux2_1 _09285_ (.A0(\top.histogram.total[18] ),
    .A1(\top.histogram.total[19] ),
    .S(net508),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05229_));
 sky130_fd_sc_hd__or2_1 _09286_ (.A(net425),
    .B(_05229_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05230_));
 sky130_fd_sc_hd__o221a_1 _09287_ (.A1(\top.histogram.total[16] ),
    .A2(net402),
    .B1(net323),
    .B2(\top.histogram.total[17] ),
    .C1(net429),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05231_));
 sky130_fd_sc_hd__a22o_1 _09288_ (.A1(net504),
    .A2(_05228_),
    .B1(_05230_),
    .B2(_05231_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05232_));
 sky130_fd_sc_hd__mux4_1 _09289_ (.A0(\top.histogram.total[28] ),
    .A1(\top.histogram.total[29] ),
    .A2(\top.histogram.total[30] ),
    .A3(\top.histogram.total[31] ),
    .S0(net509),
    .S1(net506),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05233_));
 sky130_fd_sc_hd__mux2_1 _09290_ (.A0(\top.histogram.total[26] ),
    .A1(\top.histogram.total[27] ),
    .S(net509),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05234_));
 sky130_fd_sc_hd__or2_1 _09291_ (.A(net425),
    .B(_05234_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05235_));
 sky130_fd_sc_hd__o221a_1 _09292_ (.A1(\top.histogram.total[24] ),
    .A2(net402),
    .B1(net323),
    .B2(\top.histogram.total[25] ),
    .C1(net429),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05236_));
 sky130_fd_sc_hd__a22o_1 _09293_ (.A1(net504),
    .A2(_05233_),
    .B1(_05235_),
    .B2(_05236_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05237_));
 sky130_fd_sc_hd__mux2_1 _09294_ (.A0(_05232_),
    .A1(_05237_),
    .S(net502),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05238_));
 sky130_fd_sc_hd__mux2_1 _09295_ (.A0(\top.histogram.total[2] ),
    .A1(\top.histogram.total[3] ),
    .S(net509),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05239_));
 sky130_fd_sc_hd__or2_1 _09296_ (.A(net425),
    .B(_05239_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05240_));
 sky130_fd_sc_hd__mux4_1 _09297_ (.A0(\top.histogram.total[4] ),
    .A1(\top.histogram.total[5] ),
    .A2(\top.histogram.total[6] ),
    .A3(\top.histogram.total[7] ),
    .S0(net509),
    .S1(net506),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05241_));
 sky130_fd_sc_hd__o221a_1 _09298_ (.A1(\top.histogram.total[0] ),
    .A2(net403),
    .B1(net323),
    .B2(\top.histogram.total[1] ),
    .C1(net429),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05242_));
 sky130_fd_sc_hd__a22o_1 _09299_ (.A1(net504),
    .A2(_05241_),
    .B1(_05242_),
    .B2(_05240_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05243_));
 sky130_fd_sc_hd__mux4_1 _09300_ (.A0(\top.histogram.total[8] ),
    .A1(\top.histogram.total[9] ),
    .A2(\top.histogram.total[10] ),
    .A3(\top.histogram.total[11] ),
    .S0(net509),
    .S1(net506),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05244_));
 sky130_fd_sc_hd__mux4_1 _09301_ (.A0(\top.histogram.total[12] ),
    .A1(\top.histogram.total[13] ),
    .A2(\top.histogram.total[14] ),
    .A3(\top.histogram.total[15] ),
    .S0(net509),
    .S1(net506),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05245_));
 sky130_fd_sc_hd__mux2_1 _09302_ (.A0(_05244_),
    .A1(_05245_),
    .S(net504),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05246_));
 sky130_fd_sc_hd__mux2_1 _09303_ (.A0(_05243_),
    .A1(_05246_),
    .S(net502),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05247_));
 sky130_fd_sc_hd__mux2_1 _09304_ (.A0(_05247_),
    .A1(_05238_),
    .S(\top.translation.index[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05248_));
 sky130_fd_sc_hd__a21oi_1 _09305_ (.A1(\top.translation.totalEn ),
    .A2(_05248_),
    .B1(_05227_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05249_));
 sky130_fd_sc_hd__o21ai_1 _09306_ (.A1(net513),
    .A2(_05249_),
    .B1(net423),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05250_));
 sky130_fd_sc_hd__a31o_1 _09307_ (.A1(\top.header_synthesis.bit1 ),
    .A2(net36),
    .A3(\top.header_synthesis.enable ),
    .B1(_02807_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05251_));
 sky130_fd_sc_hd__and2_1 _09308_ (.A(_05250_),
    .B(_05251_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\top.translation.writeBin ));
 sky130_fd_sc_hd__and4bb_1 _09309_ (.A_N(\top.translation.resEn ),
    .B_N(\top.translation.totalEn ),
    .C(_02807_),
    .D(_05028_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\top.controller.fin_TRN ));
 sky130_fd_sc_hd__a21bo_1 _09310_ (.A1(\top.header_synthesis.write_zeroes ),
    .A2(_05194_),
    .B1_N(_03388_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\top.header_synthesis.next_write_zeroes ));
 sky130_fd_sc_hd__and2_1 _09311_ (.A(net754),
    .B(net589),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00053_));
 sky130_fd_sc_hd__and3b_1 _09312_ (.A_N(_05052_),
    .B(_00053_),
    .C(net256),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05252_));
 sky130_fd_sc_hd__or3b_2 _09313_ (.A(_04257_),
    .B(_05052_),
    .C_N(_00053_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05253_));
 sky130_fd_sc_hd__nor2_1 _09314_ (.A(_02851_),
    .B(net220),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05254_));
 sky130_fd_sc_hd__a22o_1 _09315_ (.A1(net1002),
    .A2(net224),
    .B1(net215),
    .B2(_04515_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01248_));
 sky130_fd_sc_hd__a22o_1 _09316_ (.A1(net1096),
    .A2(net224),
    .B1(net215),
    .B2(_04511_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01249_));
 sky130_fd_sc_hd__a22o_1 _09317_ (.A1(net1109),
    .A2(net224),
    .B1(net215),
    .B2(_04507_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01250_));
 sky130_fd_sc_hd__a22o_1 _09318_ (.A1(net1027),
    .A2(net224),
    .B1(net216),
    .B2(_04503_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01251_));
 sky130_fd_sc_hd__a22o_1 _09319_ (.A1(net992),
    .A2(net224),
    .B1(net216),
    .B2(_04499_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01252_));
 sky130_fd_sc_hd__a22o_1 _09320_ (.A1(net1049),
    .A2(net224),
    .B1(net216),
    .B2(_04495_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01253_));
 sky130_fd_sc_hd__a22o_1 _09321_ (.A1(net1035),
    .A2(net224),
    .B1(net216),
    .B2(_04491_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01254_));
 sky130_fd_sc_hd__a22o_1 _09322_ (.A1(net996),
    .A2(net224),
    .B1(net216),
    .B2(_04487_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01255_));
 sky130_fd_sc_hd__a22o_1 _09323_ (.A1(net1003),
    .A2(net226),
    .B1(net217),
    .B2(_04483_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01256_));
 sky130_fd_sc_hd__a22o_1 _09324_ (.A1(net993),
    .A2(net224),
    .B1(net217),
    .B2(_04479_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01257_));
 sky130_fd_sc_hd__a22o_1 _09325_ (.A1(net995),
    .A2(net224),
    .B1(net216),
    .B2(_04475_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01258_));
 sky130_fd_sc_hd__a22o_1 _09326_ (.A1(net1017),
    .A2(net226),
    .B1(net217),
    .B2(_04471_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01259_));
 sky130_fd_sc_hd__a22o_1 _09327_ (.A1(net979),
    .A2(net226),
    .B1(net218),
    .B2(_04467_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01260_));
 sky130_fd_sc_hd__a22o_1 _09328_ (.A1(net989),
    .A2(net226),
    .B1(net217),
    .B2(_04463_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01261_));
 sky130_fd_sc_hd__a22o_1 _09329_ (.A1(net1025),
    .A2(net227),
    .B1(net218),
    .B2(_04459_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01262_));
 sky130_fd_sc_hd__a22o_1 _09330_ (.A1(net1021),
    .A2(net226),
    .B1(net217),
    .B2(_04455_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01263_));
 sky130_fd_sc_hd__a22o_1 _09331_ (.A1(net1028),
    .A2(net226),
    .B1(net218),
    .B2(_04451_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01264_));
 sky130_fd_sc_hd__a22o_1 _09332_ (.A1(net974),
    .A2(net226),
    .B1(net218),
    .B2(_04447_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01265_));
 sky130_fd_sc_hd__a22o_1 _09333_ (.A1(net1252),
    .A2(net226),
    .B1(net218),
    .B2(_04443_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01266_));
 sky130_fd_sc_hd__a22o_1 _09334_ (.A1(net1363),
    .A2(net223),
    .B1(net214),
    .B2(_04439_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01267_));
 sky130_fd_sc_hd__a22o_1 _09335_ (.A1(net1415),
    .A2(net223),
    .B1(net214),
    .B2(_04435_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01268_));
 sky130_fd_sc_hd__a22o_1 _09336_ (.A1(net998),
    .A2(net221),
    .B1(net219),
    .B2(_04431_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01269_));
 sky130_fd_sc_hd__a22o_1 _09337_ (.A1(net987),
    .A2(net222),
    .B1(net219),
    .B2(_04427_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01270_));
 sky130_fd_sc_hd__a22o_1 _09338_ (.A1(net1006),
    .A2(net221),
    .B1(net214),
    .B2(_04423_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01271_));
 sky130_fd_sc_hd__a22o_1 _09339_ (.A1(net1516),
    .A2(net223),
    .B1(net214),
    .B2(_04419_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01272_));
 sky130_fd_sc_hd__a22o_1 _09340_ (.A1(net983),
    .A2(net221),
    .B1(net219),
    .B2(_04415_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01273_));
 sky130_fd_sc_hd__a22o_1 _09341_ (.A1(net986),
    .A2(net220),
    .B1(net214),
    .B2(_04411_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01274_));
 sky130_fd_sc_hd__a22o_1 _09342_ (.A1(net964),
    .A2(net220),
    .B1(net214),
    .B2(_04407_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01275_));
 sky130_fd_sc_hd__a22o_1 _09343_ (.A1(net1629),
    .A2(net220),
    .B1(net214),
    .B2(_04403_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01276_));
 sky130_fd_sc_hd__a22o_1 _09344_ (.A1(net1795),
    .A2(net220),
    .B1(net214),
    .B2(_04399_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01277_));
 sky130_fd_sc_hd__a22o_1 _09345_ (.A1(\top.hTree.node_reg[30] ),
    .A2(net220),
    .B1(net214),
    .B2(_04395_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01278_));
 sky130_fd_sc_hd__a22o_1 _09346_ (.A1(\top.hTree.node_reg[31] ),
    .A2(net220),
    .B1(net214),
    .B2(_04391_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01279_));
 sky130_fd_sc_hd__a22o_1 _09347_ (.A1(net973),
    .A2(net225),
    .B1(net215),
    .B2(_04387_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01280_));
 sky130_fd_sc_hd__a22o_1 _09348_ (.A1(net1001),
    .A2(net225),
    .B1(net215),
    .B2(_04383_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01281_));
 sky130_fd_sc_hd__a22o_1 _09349_ (.A1(net1016),
    .A2(net225),
    .B1(net215),
    .B2(_04379_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01282_));
 sky130_fd_sc_hd__a22o_1 _09350_ (.A1(net976),
    .A2(net225),
    .B1(net215),
    .B2(_04375_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01283_));
 sky130_fd_sc_hd__a22o_1 _09351_ (.A1(net1020),
    .A2(net225),
    .B1(net215),
    .B2(_04371_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01284_));
 sky130_fd_sc_hd__a22o_1 _09352_ (.A1(net1288),
    .A2(net225),
    .B1(net215),
    .B2(_04367_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01285_));
 sky130_fd_sc_hd__a22o_1 _09353_ (.A1(net1475),
    .A2(net225),
    .B1(net215),
    .B2(_04363_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01286_));
 sky130_fd_sc_hd__a22o_1 _09354_ (.A1(net1007),
    .A2(net227),
    .B1(net216),
    .B2(_04359_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01287_));
 sky130_fd_sc_hd__a22o_1 _09355_ (.A1(net1014),
    .A2(net227),
    .B1(net217),
    .B2(_04355_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01288_));
 sky130_fd_sc_hd__a22o_1 _09356_ (.A1(net1008),
    .A2(net225),
    .B1(net217),
    .B2(_04351_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01289_));
 sky130_fd_sc_hd__a22o_1 _09357_ (.A1(net1015),
    .A2(net225),
    .B1(net217),
    .B2(_04347_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01290_));
 sky130_fd_sc_hd__a22o_1 _09358_ (.A1(net984),
    .A2(net227),
    .B1(net217),
    .B2(_04343_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01291_));
 sky130_fd_sc_hd__a22o_1 _09359_ (.A1(net982),
    .A2(net226),
    .B1(net217),
    .B2(_04339_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01292_));
 sky130_fd_sc_hd__a22o_1 _09360_ (.A1(net969),
    .A2(net226),
    .B1(net218),
    .B2(_04334_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01293_));
 sky130_fd_sc_hd__mux2_1 _09361_ (.A0(\top.hTree.nulls[46] ),
    .A1(_04331_),
    .S(net398),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05255_));
 sky130_fd_sc_hd__mux2_1 _09362_ (.A0(net1488),
    .A1(_05255_),
    .S(net228),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02298_));
 sky130_fd_sc_hd__nand2_1 _09363_ (.A(net401),
    .B(_04327_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05256_));
 sky130_fd_sc_hd__o21a_1 _09364_ (.A1(\top.hTree.nulls[47] ),
    .A2(net401),
    .B1(net229),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05257_));
 sky130_fd_sc_hd__a22o_1 _09365_ (.A1(net1665),
    .A2(net221),
    .B1(_05256_),
    .B2(_05257_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02299_));
 sky130_fd_sc_hd__nand2_1 _09366_ (.A(net398),
    .B(_04322_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05258_));
 sky130_fd_sc_hd__o21a_1 _09367_ (.A1(\top.hTree.nulls[48] ),
    .A2(net398),
    .B1(net229),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05259_));
 sky130_fd_sc_hd__a22o_1 _09368_ (.A1(net1405),
    .A2(net222),
    .B1(_05258_),
    .B2(_05259_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02300_));
 sky130_fd_sc_hd__nand2_1 _09369_ (.A(net398),
    .B(_04317_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05260_));
 sky130_fd_sc_hd__o21a_1 _09370_ (.A1(\top.hTree.nulls[49] ),
    .A2(net398),
    .B1(net228),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05261_));
 sky130_fd_sc_hd__a22o_1 _09371_ (.A1(net1275),
    .A2(net222),
    .B1(_05260_),
    .B2(_05261_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02301_));
 sky130_fd_sc_hd__nand2_1 _09372_ (.A(net398),
    .B(_04312_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05262_));
 sky130_fd_sc_hd__o21a_1 _09373_ (.A1(\top.hTree.nulls[50] ),
    .A2(net398),
    .B1(net229),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05263_));
 sky130_fd_sc_hd__a22o_1 _09374_ (.A1(net1038),
    .A2(net222),
    .B1(_05262_),
    .B2(_05263_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02302_));
 sky130_fd_sc_hd__nand2_1 _09375_ (.A(net398),
    .B(_04307_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05264_));
 sky130_fd_sc_hd__o21a_1 _09376_ (.A1(\top.hTree.nulls[51] ),
    .A2(net399),
    .B1(net228),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05265_));
 sky130_fd_sc_hd__a22o_1 _09377_ (.A1(net1030),
    .A2(net221),
    .B1(_05264_),
    .B2(_05265_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02303_));
 sky130_fd_sc_hd__nand2_1 _09378_ (.A(net398),
    .B(_04302_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05266_));
 sky130_fd_sc_hd__o21a_1 _09379_ (.A1(\top.hTree.nulls[52] ),
    .A2(net399),
    .B1(net228),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05267_));
 sky130_fd_sc_hd__a22o_1 _09380_ (.A1(net1022),
    .A2(net222),
    .B1(_05266_),
    .B2(_05267_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02304_));
 sky130_fd_sc_hd__mux2_1 _09381_ (.A0(\top.hTree.nulls[53] ),
    .A1(_04298_),
    .S(net400),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05268_));
 sky130_fd_sc_hd__mux2_1 _09382_ (.A0(net960),
    .A1(_05268_),
    .S(net228),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02305_));
 sky130_fd_sc_hd__o221a_1 _09383_ (.A1(\top.findLeastValue.least2[8] ),
    .A2(net390),
    .B1(net265),
    .B2(\top.hTree.tree_reg[54] ),
    .C1(net401),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05269_));
 sky130_fd_sc_hd__a211o_1 _09384_ (.A1(net1212),
    .A2(_02851_),
    .B1(net220),
    .C1(_05269_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05270_));
 sky130_fd_sc_hd__o21a_1 _09385_ (.A1(net1244),
    .A2(net228),
    .B1(_05270_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02306_));
 sky130_fd_sc_hd__nand2_1 _09386_ (.A(net399),
    .B(_04292_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05271_));
 sky130_fd_sc_hd__o21a_1 _09387_ (.A1(\top.hTree.nulls[55] ),
    .A2(net398),
    .B1(net228),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05272_));
 sky130_fd_sc_hd__a22o_1 _09388_ (.A1(net1024),
    .A2(net221),
    .B1(_05271_),
    .B2(_05272_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02307_));
 sky130_fd_sc_hd__nand2_1 _09389_ (.A(net399),
    .B(_04287_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05273_));
 sky130_fd_sc_hd__o21a_1 _09390_ (.A1(\top.hTree.nulls[56] ),
    .A2(net399),
    .B1(net228),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05274_));
 sky130_fd_sc_hd__a22o_1 _09391_ (.A1(net1019),
    .A2(net221),
    .B1(_05273_),
    .B2(_05274_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02308_));
 sky130_fd_sc_hd__nand2_1 _09392_ (.A(net399),
    .B(_04282_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05275_));
 sky130_fd_sc_hd__o21a_1 _09393_ (.A1(\top.hTree.nulls[57] ),
    .A2(net399),
    .B1(net229),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05276_));
 sky130_fd_sc_hd__a22o_1 _09394_ (.A1(net978),
    .A2(net221),
    .B1(_05275_),
    .B2(_05276_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02309_));
 sky130_fd_sc_hd__nand2_1 _09395_ (.A(net400),
    .B(_04277_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05277_));
 sky130_fd_sc_hd__o21a_1 _09396_ (.A1(\top.hTree.nulls[58] ),
    .A2(net400),
    .B1(net228),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05278_));
 sky130_fd_sc_hd__a22o_1 _09397_ (.A1(net990),
    .A2(net221),
    .B1(_05277_),
    .B2(_05278_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02310_));
 sky130_fd_sc_hd__nand2_1 _09398_ (.A(net400),
    .B(_04272_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05279_));
 sky130_fd_sc_hd__o21a_1 _09399_ (.A1(\top.hTree.nulls[59] ),
    .A2(net400),
    .B1(net228),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05280_));
 sky130_fd_sc_hd__a22o_1 _09400_ (.A1(net975),
    .A2(net220),
    .B1(_05279_),
    .B2(_05280_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02311_));
 sky130_fd_sc_hd__nand2_1 _09401_ (.A(net401),
    .B(_04267_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05281_));
 sky130_fd_sc_hd__o21a_1 _09402_ (.A1(\top.hTree.nulls[60] ),
    .A2(net401),
    .B1(net229),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05282_));
 sky130_fd_sc_hd__a22o_1 _09403_ (.A1(net1029),
    .A2(net221),
    .B1(_05281_),
    .B2(_05282_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02312_));
 sky130_fd_sc_hd__mux2_1 _09404_ (.A0(\top.hTree.nulls[61] ),
    .A1(_04263_),
    .S(net401),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05283_));
 sky130_fd_sc_hd__mux2_1 _09405_ (.A0(net999),
    .A1(_05283_),
    .S(net229),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02313_));
 sky130_fd_sc_hd__mux2_1 _09406_ (.A0(\top.hTree.nulls[62] ),
    .A1(_04260_),
    .S(net401),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05284_));
 sky130_fd_sc_hd__mux2_1 _09407_ (.A0(net988),
    .A1(_05284_),
    .S(net229),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02314_));
 sky130_fd_sc_hd__nor2_1 _09408_ (.A(_02851_),
    .B(_04252_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05285_));
 sky130_fd_sc_hd__a211o_1 _09409_ (.A1(\top.hTree.nulls[63] ),
    .A2(_02851_),
    .B1(net220),
    .C1(_05285_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_05286_));
 sky130_fd_sc_hd__o21a_1 _09410_ (.A1(net1580),
    .A2(net229),
    .B1(_05286_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02315_));
 sky130_fd_sc_hd__clkbuf_1 _09411_ (.A(net961),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02181_));
 sky130_fd_sc_hd__clkbuf_1 _09412_ (.A(net958),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02180_));
 sky130_fd_sc_hd__clkbuf_1 _09413_ (.A(net968),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02179_));
 sky130_fd_sc_hd__clkbuf_1 _09414_ (.A(net971),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02178_));
 sky130_fd_sc_hd__clkbuf_1 _09415_ (.A(net967),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02177_));
 sky130_fd_sc_hd__clkbuf_1 _09416_ (.A(net970),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02176_));
 sky130_fd_sc_hd__clkbuf_1 _09417_ (.A(net972),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02175_));
 sky130_fd_sc_hd__clkbuf_1 _09418_ (.A(net962),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02174_));
 sky130_fd_sc_hd__clkbuf_1 _09419_ (.A(net965),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02173_));
 sky130_fd_sc_hd__clkbuf_1 _09420_ (.A(net963),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02172_));
 sky130_fd_sc_hd__clkbuf_1 _09421_ (.A(net959),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02171_));
 sky130_fd_sc_hd__clkbuf_1 _09422_ (.A(net966),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_02170_));
 sky130_fd_sc_hd__and2_1 _09423_ (.A(net754),
    .B(net589),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00054_));
 sky130_fd_sc_hd__and2_1 _09424_ (.A(net747),
    .B(net582),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00055_));
 sky130_fd_sc_hd__and2_1 _09425_ (.A(net754),
    .B(net589),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00056_));
 sky130_fd_sc_hd__and2_1 _09426_ (.A(net747),
    .B(net582),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00057_));
 sky130_fd_sc_hd__and2_1 _09427_ (.A(net747),
    .B(net582),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00058_));
 sky130_fd_sc_hd__and2_1 _09428_ (.A(net801),
    .B(net636),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00059_));
 sky130_fd_sc_hd__and2_1 _09429_ (.A(net801),
    .B(net636),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00060_));
 sky130_fd_sc_hd__and2_1 _09430_ (.A(net755),
    .B(net590),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00061_));
 sky130_fd_sc_hd__and2_1 _09431_ (.A(net755),
    .B(net590),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00062_));
 sky130_fd_sc_hd__and2_1 _09432_ (.A(net746),
    .B(net581),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00063_));
 sky130_fd_sc_hd__and2_1 _09433_ (.A(net746),
    .B(net581),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00064_));
 sky130_fd_sc_hd__and2_1 _09434_ (.A(net746),
    .B(net581),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00065_));
 sky130_fd_sc_hd__and2_1 _09435_ (.A(net751),
    .B(net586),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00066_));
 sky130_fd_sc_hd__and2_1 _09436_ (.A(net741),
    .B(net576),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00067_));
 sky130_fd_sc_hd__and2_1 _09437_ (.A(net741),
    .B(net576),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00068_));
 sky130_fd_sc_hd__and2_1 _09438_ (.A(net733),
    .B(net568),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00069_));
 sky130_fd_sc_hd__and2_1 _09439_ (.A(net724),
    .B(net559),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00070_));
 sky130_fd_sc_hd__and2_1 _09440_ (.A(net724),
    .B(net559),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00071_));
 sky130_fd_sc_hd__and2_1 _09441_ (.A(net724),
    .B(net559),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00072_));
 sky130_fd_sc_hd__and2_1 _09442_ (.A(net724),
    .B(net559),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00073_));
 sky130_fd_sc_hd__and2_1 _09443_ (.A(net726),
    .B(net561),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00074_));
 sky130_fd_sc_hd__and2_1 _09444_ (.A(net742),
    .B(net577),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00075_));
 sky130_fd_sc_hd__and2_1 _09445_ (.A(net742),
    .B(net577),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00076_));
 sky130_fd_sc_hd__and2_1 _09446_ (.A(net750),
    .B(net585),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00077_));
 sky130_fd_sc_hd__and2_1 _09447_ (.A(net750),
    .B(net585),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00078_));
 sky130_fd_sc_hd__and2_1 _09448_ (.A(net750),
    .B(net585),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00079_));
 sky130_fd_sc_hd__and2_1 _09449_ (.A(net750),
    .B(net585),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00080_));
 sky130_fd_sc_hd__and2_1 _09450_ (.A(net741),
    .B(net576),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00081_));
 sky130_fd_sc_hd__and2_1 _09451_ (.A(net741),
    .B(net576),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00082_));
 sky130_fd_sc_hd__and2_1 _09452_ (.A(net751),
    .B(net586),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00083_));
 sky130_fd_sc_hd__and2_1 _09453_ (.A(net751),
    .B(net586),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00084_));
 sky130_fd_sc_hd__and2_1 _09454_ (.A(net732),
    .B(net567),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00085_));
 sky130_fd_sc_hd__and2_1 _09455_ (.A(net758),
    .B(net593),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00086_));
 sky130_fd_sc_hd__and2_1 _09456_ (.A(net730),
    .B(net565),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00087_));
 sky130_fd_sc_hd__and2_1 _09457_ (.A(net730),
    .B(net565),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00088_));
 sky130_fd_sc_hd__and2_1 _09458_ (.A(net731),
    .B(net566),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00089_));
 sky130_fd_sc_hd__and2_1 _09459_ (.A(net731),
    .B(net566),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00090_));
 sky130_fd_sc_hd__and2_1 _09460_ (.A(net732),
    .B(net567),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00091_));
 sky130_fd_sc_hd__and2_1 _09461_ (.A(net842),
    .B(net677),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00092_));
 sky130_fd_sc_hd__and2_1 _09462_ (.A(net838),
    .B(net673),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00093_));
 sky130_fd_sc_hd__and2_1 _09463_ (.A(net836),
    .B(net671),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00094_));
 sky130_fd_sc_hd__and2_1 _09464_ (.A(net840),
    .B(net675),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00095_));
 sky130_fd_sc_hd__and2_1 _09465_ (.A(net842),
    .B(net677),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00096_));
 sky130_fd_sc_hd__and2_1 _09466_ (.A(net842),
    .B(net677),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00097_));
 sky130_fd_sc_hd__and2_1 _09467_ (.A(net842),
    .B(net677),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00098_));
 sky130_fd_sc_hd__and2_1 _09468_ (.A(net840),
    .B(net675),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00099_));
 sky130_fd_sc_hd__and2_1 _09469_ (.A(net811),
    .B(net646),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00100_));
 sky130_fd_sc_hd__and2_1 _09470_ (.A(net837),
    .B(net672),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00101_));
 sky130_fd_sc_hd__and2_1 _09471_ (.A(net838),
    .B(net673),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00102_));
 sky130_fd_sc_hd__and2_1 _09472_ (.A(net837),
    .B(net672),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00103_));
 sky130_fd_sc_hd__and2_1 _09473_ (.A(net837),
    .B(net672),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00104_));
 sky130_fd_sc_hd__and2_1 _09474_ (.A(net811),
    .B(net646),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00105_));
 sky130_fd_sc_hd__and2_1 _09475_ (.A(net785),
    .B(net620),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00106_));
 sky130_fd_sc_hd__and2_1 _09476_ (.A(net785),
    .B(net620),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00107_));
 sky130_fd_sc_hd__and2_1 _09477_ (.A(net784),
    .B(net619),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00108_));
 sky130_fd_sc_hd__and2_1 _09478_ (.A(net811),
    .B(net646),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00109_));
 sky130_fd_sc_hd__and2_1 _09479_ (.A(net778),
    .B(net613),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00110_));
 sky130_fd_sc_hd__and2_1 _09480_ (.A(net779),
    .B(net614),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00111_));
 sky130_fd_sc_hd__and2_1 _09481_ (.A(net765),
    .B(net600),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00112_));
 sky130_fd_sc_hd__and2_1 _09482_ (.A(net778),
    .B(net613),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00113_));
 sky130_fd_sc_hd__and2_1 _09483_ (.A(net765),
    .B(net600),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00114_));
 sky130_fd_sc_hd__and2_1 _09484_ (.A(net765),
    .B(net600),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00115_));
 sky130_fd_sc_hd__and2_1 _09485_ (.A(net778),
    .B(net613),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00116_));
 sky130_fd_sc_hd__and2_1 _09486_ (.A(net765),
    .B(net600),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00117_));
 sky130_fd_sc_hd__and2_1 _09487_ (.A(net778),
    .B(net613),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00118_));
 sky130_fd_sc_hd__and2_1 _09488_ (.A(net778),
    .B(net613),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00119_));
 sky130_fd_sc_hd__and2_1 _09489_ (.A(net778),
    .B(net613),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00120_));
 sky130_fd_sc_hd__and2_1 _09490_ (.A(net778),
    .B(net613),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00121_));
 sky130_fd_sc_hd__and2_1 _09491_ (.A(net765),
    .B(net600),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00122_));
 sky130_fd_sc_hd__and2_1 _09492_ (.A(net778),
    .B(net613),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00123_));
 sky130_fd_sc_hd__and2_1 _09493_ (.A(net780),
    .B(net615),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00124_));
 sky130_fd_sc_hd__and2_1 _09494_ (.A(net780),
    .B(net615),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00125_));
 sky130_fd_sc_hd__and2_1 _09495_ (.A(net779),
    .B(net614),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00126_));
 sky130_fd_sc_hd__and2_1 _09496_ (.A(net779),
    .B(net614),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00127_));
 sky130_fd_sc_hd__and2_1 _09497_ (.A(net727),
    .B(net562),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00128_));
 sky130_fd_sc_hd__and2_1 _09498_ (.A(net729),
    .B(net564),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00129_));
 sky130_fd_sc_hd__and2_1 _09499_ (.A(net729),
    .B(net564),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00130_));
 sky130_fd_sc_hd__and2_1 _09500_ (.A(net729),
    .B(net564),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00131_));
 sky130_fd_sc_hd__and2_1 _09501_ (.A(net729),
    .B(net564),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00132_));
 sky130_fd_sc_hd__and2_1 _09502_ (.A(net727),
    .B(net562),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00133_));
 sky130_fd_sc_hd__and2_1 _09503_ (.A(net730),
    .B(net565),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00134_));
 sky130_fd_sc_hd__and2_1 _09504_ (.A(net728),
    .B(net563),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00135_));
 sky130_fd_sc_hd__and2_1 _09505_ (.A(net732),
    .B(net567),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00136_));
 sky130_fd_sc_hd__and2_1 _09506_ (.A(net732),
    .B(net567),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00137_));
 sky130_fd_sc_hd__and2_1 _09507_ (.A(net752),
    .B(net587),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00138_));
 sky130_fd_sc_hd__and2_1 _09508_ (.A(net733),
    .B(net568),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00139_));
 sky130_fd_sc_hd__and2_1 _09509_ (.A(net752),
    .B(net587),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00140_));
 sky130_fd_sc_hd__and2_1 _09510_ (.A(net735),
    .B(net570),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00141_));
 sky130_fd_sc_hd__and2_1 _09511_ (.A(net732),
    .B(net567),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00142_));
 sky130_fd_sc_hd__and2_1 _09512_ (.A(net752),
    .B(net587),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00143_));
 sky130_fd_sc_hd__and2_1 _09513_ (.A(net732),
    .B(net567),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00144_));
 sky130_fd_sc_hd__and2_1 _09514_ (.A(net734),
    .B(net569),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00145_));
 sky130_fd_sc_hd__and2_1 _09515_ (.A(net733),
    .B(net568),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00146_));
 sky130_fd_sc_hd__and2_1 _09516_ (.A(net735),
    .B(net570),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00147_));
 sky130_fd_sc_hd__and2_1 _09517_ (.A(net752),
    .B(net587),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00148_));
 sky130_fd_sc_hd__and2_1 _09518_ (.A(net734),
    .B(net569),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00149_));
 sky130_fd_sc_hd__and2_1 _09519_ (.A(net752),
    .B(net587),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00150_));
 sky130_fd_sc_hd__and2_1 _09520_ (.A(net735),
    .B(net570),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00151_));
 sky130_fd_sc_hd__and2_1 _09521_ (.A(net752),
    .B(net587),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00152_));
 sky130_fd_sc_hd__and2_1 _09522_ (.A(net745),
    .B(net580),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00153_));
 sky130_fd_sc_hd__and2_1 _09523_ (.A(net743),
    .B(net578),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00154_));
 sky130_fd_sc_hd__and2_1 _09524_ (.A(net797),
    .B(net632),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00155_));
 sky130_fd_sc_hd__and2_1 _09525_ (.A(net745),
    .B(net580),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00156_));
 sky130_fd_sc_hd__and2_1 _09526_ (.A(net747),
    .B(net582),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00157_));
 sky130_fd_sc_hd__and2_1 _09527_ (.A(net747),
    .B(net582),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00158_));
 sky130_fd_sc_hd__and2_1 _09528_ (.A(net797),
    .B(net632),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00159_));
 sky130_fd_sc_hd__and2_1 _09529_ (.A(net801),
    .B(net636),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00160_));
 sky130_fd_sc_hd__and2_1 _09530_ (.A(net744),
    .B(net579),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00161_));
 sky130_fd_sc_hd__and2_1 _09531_ (.A(net743),
    .B(net578),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00162_));
 sky130_fd_sc_hd__and2_1 _09532_ (.A(net744),
    .B(net579),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00163_));
 sky130_fd_sc_hd__and2_1 _09533_ (.A(net744),
    .B(net579),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00164_));
 sky130_fd_sc_hd__and2_1 _09534_ (.A(net746),
    .B(net581),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00165_));
 sky130_fd_sc_hd__and2_1 _09535_ (.A(net741),
    .B(net576),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00166_));
 sky130_fd_sc_hd__and2_1 _09536_ (.A(net744),
    .B(net579),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00167_));
 sky130_fd_sc_hd__and2_1 _09537_ (.A(net744),
    .B(net579),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00168_));
 sky130_fd_sc_hd__and2_1 _09538_ (.A(net737),
    .B(net572),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00169_));
 sky130_fd_sc_hd__and2_1 _09539_ (.A(net722),
    .B(net557),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00170_));
 sky130_fd_sc_hd__and2_1 _09540_ (.A(net722),
    .B(net557),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00171_));
 sky130_fd_sc_hd__and2_1 _09541_ (.A(net722),
    .B(net557),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00172_));
 sky130_fd_sc_hd__and2_1 _09542_ (.A(net722),
    .B(net557),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00173_));
 sky130_fd_sc_hd__and2_1 _09543_ (.A(net722),
    .B(net557),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00174_));
 sky130_fd_sc_hd__and2_1 _09544_ (.A(net737),
    .B(net572),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00175_));
 sky130_fd_sc_hd__and2_1 _09545_ (.A(net737),
    .B(net572),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00176_));
 sky130_fd_sc_hd__and2_1 _09546_ (.A(net737),
    .B(net572),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00177_));
 sky130_fd_sc_hd__and2_1 _09547_ (.A(net722),
    .B(net557),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00178_));
 sky130_fd_sc_hd__and2_1 _09548_ (.A(net722),
    .B(net557),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00179_));
 sky130_fd_sc_hd__and2_1 _09549_ (.A(net723),
    .B(net558),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00180_));
 sky130_fd_sc_hd__and2_1 _09550_ (.A(net737),
    .B(net572),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00181_));
 sky130_fd_sc_hd__and2_1 _09551_ (.A(net737),
    .B(net572),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00182_));
 sky130_fd_sc_hd__and2_1 _09552_ (.A(net738),
    .B(net573),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00183_));
 sky130_fd_sc_hd__and2_1 _09553_ (.A(net738),
    .B(net573),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00184_));
 sky130_fd_sc_hd__and2_1 _09554_ (.A(net729),
    .B(net564),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00185_));
 sky130_fd_sc_hd__and2_1 _09555_ (.A(net734),
    .B(net569),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00186_));
 sky130_fd_sc_hd__and2_1 _09556_ (.A(net734),
    .B(net569),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00187_));
 sky130_fd_sc_hd__and2_1 _09557_ (.A(net763),
    .B(net598),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00188_));
 sky130_fd_sc_hd__and2_1 _09558_ (.A(net763),
    .B(net598),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00189_));
 sky130_fd_sc_hd__and2_1 _09559_ (.A(net763),
    .B(net598),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00190_));
 sky130_fd_sc_hd__and2_1 _09560_ (.A(net763),
    .B(net598),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00191_));
 sky130_fd_sc_hd__and2_1 _09561_ (.A(net763),
    .B(net598),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00192_));
 sky130_fd_sc_hd__and2_1 _09562_ (.A(net763),
    .B(net598),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00193_));
 sky130_fd_sc_hd__and2_1 _09563_ (.A(net763),
    .B(net598),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00194_));
 sky130_fd_sc_hd__and2_1 _09564_ (.A(net772),
    .B(net607),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00195_));
 sky130_fd_sc_hd__and2_1 _09565_ (.A(net780),
    .B(net615),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00196_));
 sky130_fd_sc_hd__and2_1 _09566_ (.A(net774),
    .B(net609),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00197_));
 sky130_fd_sc_hd__and2_1 _09567_ (.A(net772),
    .B(net607),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00198_));
 sky130_fd_sc_hd__and2_1 _09568_ (.A(net773),
    .B(net608),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00199_));
 sky130_fd_sc_hd__and2_1 _09569_ (.A(net787),
    .B(net622),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00200_));
 sky130_fd_sc_hd__and2_1 _09570_ (.A(net788),
    .B(net623),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00201_));
 sky130_fd_sc_hd__and2_1 _09571_ (.A(net772),
    .B(net607),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00202_));
 sky130_fd_sc_hd__and2_1 _09572_ (.A(net772),
    .B(net607),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00203_));
 sky130_fd_sc_hd__and2_1 _09573_ (.A(net747),
    .B(net582),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00204_));
 sky130_fd_sc_hd__and2_1 _09574_ (.A(net747),
    .B(net582),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00205_));
 sky130_fd_sc_hd__and2_1 _09575_ (.A(net799),
    .B(net634),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00206_));
 sky130_fd_sc_hd__and2_1 _09576_ (.A(net798),
    .B(net633),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00207_));
 sky130_fd_sc_hd__and2_1 _09577_ (.A(net800),
    .B(net635),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00208_));
 sky130_fd_sc_hd__and2_1 _09578_ (.A(net798),
    .B(net633),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00209_));
 sky130_fd_sc_hd__and2_1 _09579_ (.A(net798),
    .B(net633),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00210_));
 sky130_fd_sc_hd__and2_1 _09580_ (.A(net798),
    .B(net633),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00211_));
 sky130_fd_sc_hd__and2_1 _09581_ (.A(net745),
    .B(net580),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00212_));
 sky130_fd_sc_hd__and2_1 _09582_ (.A(net748),
    .B(net583),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00213_));
 sky130_fd_sc_hd__and2_1 _09583_ (.A(net797),
    .B(net632),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00214_));
 sky130_fd_sc_hd__and2_1 _09584_ (.A(net797),
    .B(net632),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00215_));
 sky130_fd_sc_hd__and2_1 _09585_ (.A(net745),
    .B(net580),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00216_));
 sky130_fd_sc_hd__and2_1 _09586_ (.A(net743),
    .B(net578),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00217_));
 sky130_fd_sc_hd__and2_1 _09587_ (.A(net799),
    .B(net634),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00218_));
 sky130_fd_sc_hd__and2_1 _09588_ (.A(net798),
    .B(net633),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00219_));
 sky130_fd_sc_hd__and2_1 _09589_ (.A(net724),
    .B(net559),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00220_));
 sky130_fd_sc_hd__and2_1 _09590_ (.A(net724),
    .B(net559),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00221_));
 sky130_fd_sc_hd__and2_1 _09591_ (.A(net723),
    .B(net558),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00222_));
 sky130_fd_sc_hd__and2_1 _09592_ (.A(net723),
    .B(net558),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00223_));
 sky130_fd_sc_hd__and2_1 _09593_ (.A(net742),
    .B(net577),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00224_));
 sky130_fd_sc_hd__and2_1 _09594_ (.A(net726),
    .B(net561),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00225_));
 sky130_fd_sc_hd__and2_1 _09595_ (.A(net742),
    .B(net577),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00226_));
 sky130_fd_sc_hd__and2_1 _09596_ (.A(net742),
    .B(net577),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00227_));
 sky130_fd_sc_hd__and2_1 _09597_ (.A(net742),
    .B(net577),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00228_));
 sky130_fd_sc_hd__and2_1 _09598_ (.A(net742),
    .B(net577),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00229_));
 sky130_fd_sc_hd__and2_1 _09599_ (.A(net724),
    .B(net559),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00230_));
 sky130_fd_sc_hd__and2_1 _09600_ (.A(net724),
    .B(net559),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00231_));
 sky130_fd_sc_hd__and2_1 _09601_ (.A(net741),
    .B(net576),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00232_));
 sky130_fd_sc_hd__and2_1 _09602_ (.A(net741),
    .B(net576),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00233_));
 sky130_fd_sc_hd__and2_1 _09603_ (.A(net741),
    .B(net576),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00234_));
 sky130_fd_sc_hd__and2_1 _09604_ (.A(net749),
    .B(net584),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00235_));
 sky130_fd_sc_hd__and2_1 _09605_ (.A(net725),
    .B(net560),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00236_));
 sky130_fd_sc_hd__and2_1 _09606_ (.A(net725),
    .B(net560),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00237_));
 sky130_fd_sc_hd__and2_1 _09607_ (.A(net721),
    .B(net556),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00238_));
 sky130_fd_sc_hd__and2_1 _09608_ (.A(net721),
    .B(net556),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00239_));
 sky130_fd_sc_hd__and2_1 _09609_ (.A(net725),
    .B(net560),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00240_));
 sky130_fd_sc_hd__and2_1 _09610_ (.A(net725),
    .B(net560),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00241_));
 sky130_fd_sc_hd__and2_1 _09611_ (.A(net725),
    .B(net560),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00242_));
 sky130_fd_sc_hd__and2_1 _09612_ (.A(net724),
    .B(net559),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00243_));
 sky130_fd_sc_hd__and2_1 _09613_ (.A(net724),
    .B(net559),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00244_));
 sky130_fd_sc_hd__and2_1 _09614_ (.A(net726),
    .B(net561),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00245_));
 sky130_fd_sc_hd__and2_1 _09615_ (.A(net733),
    .B(net568),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00246_));
 sky130_fd_sc_hd__and2_1 _09616_ (.A(net750),
    .B(net585),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00247_));
 sky130_fd_sc_hd__and2_1 _09617_ (.A(net733),
    .B(net568),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00248_));
 sky130_fd_sc_hd__and2_1 _09618_ (.A(net769),
    .B(net604),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00249_));
 sky130_fd_sc_hd__and2_1 _09619_ (.A(net770),
    .B(net605),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00250_));
 sky130_fd_sc_hd__and2_1 _09620_ (.A(net770),
    .B(net605),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00251_));
 sky130_fd_sc_hd__and2_1 _09621_ (.A(net770),
    .B(net605),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00252_));
 sky130_fd_sc_hd__and2_1 _09622_ (.A(net769),
    .B(net604),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00253_));
 sky130_fd_sc_hd__and2_1 _09623_ (.A(net769),
    .B(net604),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00254_));
 sky130_fd_sc_hd__and2_1 _09624_ (.A(net770),
    .B(net605),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00255_));
 sky130_fd_sc_hd__and2_1 _09625_ (.A(net770),
    .B(net605),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00256_));
 sky130_fd_sc_hd__and2_1 _09626_ (.A(net756),
    .B(net591),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00257_));
 sky130_fd_sc_hd__and2_1 _09627_ (.A(net772),
    .B(net607),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00258_));
 sky130_fd_sc_hd__and2_1 _09628_ (.A(net768),
    .B(net603),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00259_));
 sky130_fd_sc_hd__and2_1 _09629_ (.A(net767),
    .B(net602),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00260_));
 sky130_fd_sc_hd__and2_1 _09630_ (.A(net767),
    .B(net602),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00261_));
 sky130_fd_sc_hd__and2_1 _09631_ (.A(net767),
    .B(net602),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00262_));
 sky130_fd_sc_hd__and2_1 _09632_ (.A(net767),
    .B(net602),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00263_));
 sky130_fd_sc_hd__and2_1 _09633_ (.A(net760),
    .B(net595),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00264_));
 sky130_fd_sc_hd__and2_1 _09634_ (.A(net760),
    .B(net595),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00265_));
 sky130_fd_sc_hd__and2_1 _09635_ (.A(net760),
    .B(net595),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00266_));
 sky130_fd_sc_hd__and2_1 _09636_ (.A(net772),
    .B(net607),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00267_));
 sky130_fd_sc_hd__and2_1 _09637_ (.A(net761),
    .B(net596),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00268_));
 sky130_fd_sc_hd__and2_1 _09638_ (.A(net761),
    .B(net596),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00269_));
 sky130_fd_sc_hd__and2_1 _09639_ (.A(net760),
    .B(net595),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00270_));
 sky130_fd_sc_hd__and2_1 _09640_ (.A(net760),
    .B(net595),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00271_));
 sky130_fd_sc_hd__and2_1 _09641_ (.A(net762),
    .B(net597),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00272_));
 sky130_fd_sc_hd__and2_1 _09642_ (.A(net761),
    .B(net596),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00273_));
 sky130_fd_sc_hd__and2_1 _09643_ (.A(net761),
    .B(net596),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00274_));
 sky130_fd_sc_hd__and2_1 _09644_ (.A(net762),
    .B(net597),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00275_));
 sky130_fd_sc_hd__and2_1 _09645_ (.A(net762),
    .B(net597),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00276_));
 sky130_fd_sc_hd__and2_1 _09646_ (.A(net768),
    .B(net603),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00277_));
 sky130_fd_sc_hd__and2_1 _09647_ (.A(net768),
    .B(net603),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00278_));
 sky130_fd_sc_hd__and2_1 _09648_ (.A(net768),
    .B(net603),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00279_));
 sky130_fd_sc_hd__and2_1 _09649_ (.A(net772),
    .B(net607),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00280_));
 sky130_fd_sc_hd__and2_1 _09650_ (.A(net787),
    .B(net622),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00281_));
 sky130_fd_sc_hd__and2_1 _09651_ (.A(net774),
    .B(net609),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00282_));
 sky130_fd_sc_hd__and2_1 _09652_ (.A(net774),
    .B(net609),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00283_));
 sky130_fd_sc_hd__and2_1 _09653_ (.A(net789),
    .B(net624),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00284_));
 sky130_fd_sc_hd__and2_1 _09654_ (.A(net774),
    .B(net609),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00285_));
 sky130_fd_sc_hd__and2_1 _09655_ (.A(net774),
    .B(net609),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00286_));
 sky130_fd_sc_hd__and2_1 _09656_ (.A(net774),
    .B(net609),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00287_));
 sky130_fd_sc_hd__and2_1 _09657_ (.A(net789),
    .B(net624),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00288_));
 sky130_fd_sc_hd__and2_1 _09658_ (.A(net787),
    .B(net622),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00289_));
 sky130_fd_sc_hd__and2_1 _09659_ (.A(net846),
    .B(net681),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00290_));
 sky130_fd_sc_hd__and2_1 _09660_ (.A(net846),
    .B(net681),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00291_));
 sky130_fd_sc_hd__and2_1 _09661_ (.A(net846),
    .B(net681),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00292_));
 sky130_fd_sc_hd__and2_1 _09662_ (.A(net848),
    .B(net683),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00293_));
 sky130_fd_sc_hd__and2_1 _09663_ (.A(net848),
    .B(net683),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00294_));
 sky130_fd_sc_hd__and2_1 _09664_ (.A(net848),
    .B(net683),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00295_));
 sky130_fd_sc_hd__and2_1 _09665_ (.A(net789),
    .B(net624),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00296_));
 sky130_fd_sc_hd__and2_1 _09666_ (.A(net788),
    .B(net623),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00297_));
 sky130_fd_sc_hd__and2_1 _09667_ (.A(net787),
    .B(net622),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00298_));
 sky130_fd_sc_hd__and2_1 _09668_ (.A(net725),
    .B(net560),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00299_));
 sky130_fd_sc_hd__and2_1 _09669_ (.A(net764),
    .B(net599),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00300_));
 sky130_fd_sc_hd__and2_1 _09670_ (.A(net733),
    .B(net568),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00301_));
 sky130_fd_sc_hd__and2_1 _09671_ (.A(net754),
    .B(net589),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00302_));
 sky130_fd_sc_hd__and2_1 _09672_ (.A(net750),
    .B(net585),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00303_));
 sky130_fd_sc_hd__and2_1 _09673_ (.A(net734),
    .B(net569),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00304_));
 sky130_fd_sc_hd__and2_1 _09674_ (.A(net727),
    .B(net562),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00305_));
 sky130_fd_sc_hd__and2_1 _09675_ (.A(net788),
    .B(net623),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00306_));
 sky130_fd_sc_hd__and2_1 _09676_ (.A(net787),
    .B(net622),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00307_));
 sky130_fd_sc_hd__and2_1 _09677_ (.A(net838),
    .B(net673),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00308_));
 sky130_fd_sc_hd__and2_1 _09678_ (.A(net850),
    .B(net685),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00309_));
 sky130_fd_sc_hd__and2_1 _09679_ (.A(net842),
    .B(net677),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00310_));
 sky130_fd_sc_hd__and2_1 _09680_ (.A(net843),
    .B(net678),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00311_));
 sky130_fd_sc_hd__and2_1 _09681_ (.A(net843),
    .B(net678),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00312_));
 sky130_fd_sc_hd__and2_1 _09682_ (.A(net843),
    .B(net678),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00313_));
 sky130_fd_sc_hd__and2_1 _09683_ (.A(net856),
    .B(net691),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00314_));
 sky130_fd_sc_hd__and2_1 _09684_ (.A(net862),
    .B(net697),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00315_));
 sky130_fd_sc_hd__and2_1 _09685_ (.A(net863),
    .B(net698),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00316_));
 sky130_fd_sc_hd__and2_1 _09686_ (.A(net870),
    .B(net705),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00317_));
 sky130_fd_sc_hd__and2_1 _09687_ (.A(net870),
    .B(net705),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00318_));
 sky130_fd_sc_hd__and2_1 _09688_ (.A(net873),
    .B(net708),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00319_));
 sky130_fd_sc_hd__and2_1 _09689_ (.A(net873),
    .B(net708),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00320_));
 sky130_fd_sc_hd__and2_1 _09690_ (.A(net874),
    .B(net709),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00321_));
 sky130_fd_sc_hd__and2_1 _09691_ (.A(net868),
    .B(net703),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00322_));
 sky130_fd_sc_hd__and2_1 _09692_ (.A(net869),
    .B(net704),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00323_));
 sky130_fd_sc_hd__and2_1 _09693_ (.A(net868),
    .B(net703),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00324_));
 sky130_fd_sc_hd__and2_1 _09694_ (.A(net868),
    .B(net703),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00325_));
 sky130_fd_sc_hd__and2_1 _09695_ (.A(net852),
    .B(net687),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00326_));
 sky130_fd_sc_hd__and2_1 _09696_ (.A(net852),
    .B(net687),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00327_));
 sky130_fd_sc_hd__and2_1 _09697_ (.A(net853),
    .B(net688),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00328_));
 sky130_fd_sc_hd__and2_1 _09698_ (.A(net853),
    .B(net688),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00329_));
 sky130_fd_sc_hd__and2_1 _09699_ (.A(net848),
    .B(net683),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00330_));
 sky130_fd_sc_hd__and2_1 _09700_ (.A(net849),
    .B(net684),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00331_));
 sky130_fd_sc_hd__and2_1 _09701_ (.A(net848),
    .B(net683),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00332_));
 sky130_fd_sc_hd__and2_1 _09702_ (.A(net792),
    .B(net627),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00333_));
 sky130_fd_sc_hd__and2_1 _09703_ (.A(net792),
    .B(net627),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00334_));
 sky130_fd_sc_hd__and2_1 _09704_ (.A(net792),
    .B(net627),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00335_));
 sky130_fd_sc_hd__and2_1 _09705_ (.A(net792),
    .B(net627),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00336_));
 sky130_fd_sc_hd__and2_1 _09706_ (.A(net791),
    .B(net626),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00337_));
 sky130_fd_sc_hd__and2_1 _09707_ (.A(net787),
    .B(net622),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00338_));
 sky130_fd_sc_hd__and2_1 _09708_ (.A(net784),
    .B(net619),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00339_));
 sky130_fd_sc_hd__and2_1 _09709_ (.A(net839),
    .B(net674),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00340_));
 sky130_fd_sc_hd__and2_1 _09710_ (.A(net842),
    .B(net677),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00341_));
 sky130_fd_sc_hd__and2_1 _09711_ (.A(net842),
    .B(net677),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00342_));
 sky130_fd_sc_hd__and2_1 _09712_ (.A(net856),
    .B(net691),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00343_));
 sky130_fd_sc_hd__and2_1 _09713_ (.A(net857),
    .B(net692),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00344_));
 sky130_fd_sc_hd__and2_1 _09714_ (.A(net864),
    .B(net699),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00345_));
 sky130_fd_sc_hd__and2_1 _09715_ (.A(net864),
    .B(net699),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00346_));
 sky130_fd_sc_hd__and2_1 _09716_ (.A(net862),
    .B(net697),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00347_));
 sky130_fd_sc_hd__and2_1 _09717_ (.A(net863),
    .B(net698),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00348_));
 sky130_fd_sc_hd__and2_1 _09718_ (.A(net872),
    .B(net707),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00349_));
 sky130_fd_sc_hd__and2_1 _09719_ (.A(net870),
    .B(net705),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00350_));
 sky130_fd_sc_hd__and2_1 _09720_ (.A(net870),
    .B(net705),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00351_));
 sky130_fd_sc_hd__and2_1 _09721_ (.A(net870),
    .B(net705),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00352_));
 sky130_fd_sc_hd__and2_1 _09722_ (.A(net872),
    .B(net707),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00353_));
 sky130_fd_sc_hd__and2_1 _09723_ (.A(net867),
    .B(net702),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00354_));
 sky130_fd_sc_hd__and2_1 _09724_ (.A(net866),
    .B(net701),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00355_));
 sky130_fd_sc_hd__and2_1 _09725_ (.A(net866),
    .B(net701),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00356_));
 sky130_fd_sc_hd__and2_1 _09726_ (.A(net866),
    .B(net701),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00357_));
 sky130_fd_sc_hd__and2_1 _09727_ (.A(net851),
    .B(net686),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00358_));
 sky130_fd_sc_hd__and2_1 _09728_ (.A(net851),
    .B(net686),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00359_));
 sky130_fd_sc_hd__and2_1 _09729_ (.A(net851),
    .B(net686),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00360_));
 sky130_fd_sc_hd__and2_1 _09730_ (.A(net850),
    .B(net685),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00361_));
 sky130_fd_sc_hd__and2_1 _09731_ (.A(net850),
    .B(net685),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00362_));
 sky130_fd_sc_hd__and2_1 _09732_ (.A(net847),
    .B(net682),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00363_));
 sky130_fd_sc_hd__and2_1 _09733_ (.A(net846),
    .B(net681),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00364_));
 sky130_fd_sc_hd__and2_1 _09734_ (.A(net790),
    .B(net625),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00365_));
 sky130_fd_sc_hd__and2_1 _09735_ (.A(net790),
    .B(net625),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00366_));
 sky130_fd_sc_hd__and2_1 _09736_ (.A(net790),
    .B(net625),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00367_));
 sky130_fd_sc_hd__and2_1 _09737_ (.A(net790),
    .B(net625),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00368_));
 sky130_fd_sc_hd__and2_1 _09738_ (.A(net791),
    .B(net626),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00369_));
 sky130_fd_sc_hd__and2_1 _09739_ (.A(net787),
    .B(net622),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00370_));
 sky130_fd_sc_hd__and2_1 _09740_ (.A(net779),
    .B(net614),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00371_));
 sky130_fd_sc_hd__and2_1 _09741_ (.A(net838),
    .B(net673),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00372_));
 sky130_fd_sc_hd__and2_1 _09742_ (.A(net842),
    .B(net677),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00373_));
 sky130_fd_sc_hd__and2_1 _09743_ (.A(net842),
    .B(net677),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00374_));
 sky130_fd_sc_hd__and2_1 _09744_ (.A(net856),
    .B(net691),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00375_));
 sky130_fd_sc_hd__and2_1 _09745_ (.A(net856),
    .B(net691),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00376_));
 sky130_fd_sc_hd__and2_1 _09746_ (.A(net856),
    .B(net691),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00377_));
 sky130_fd_sc_hd__and2_1 _09747_ (.A(net856),
    .B(net691),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00378_));
 sky130_fd_sc_hd__and2_1 _09748_ (.A(net863),
    .B(net698),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00379_));
 sky130_fd_sc_hd__and2_1 _09749_ (.A(net863),
    .B(net698),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00380_));
 sky130_fd_sc_hd__and2_1 _09750_ (.A(net872),
    .B(net707),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00381_));
 sky130_fd_sc_hd__and2_1 _09751_ (.A(net870),
    .B(net705),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00382_));
 sky130_fd_sc_hd__and2_1 _09752_ (.A(net873),
    .B(net708),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00383_));
 sky130_fd_sc_hd__and2_1 _09753_ (.A(net873),
    .B(net708),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00384_));
 sky130_fd_sc_hd__and2_1 _09754_ (.A(net874),
    .B(net709),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00385_));
 sky130_fd_sc_hd__and2_1 _09755_ (.A(net869),
    .B(net704),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00386_));
 sky130_fd_sc_hd__and2_1 _09756_ (.A(net869),
    .B(net704),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00387_));
 sky130_fd_sc_hd__and2_1 _09757_ (.A(net868),
    .B(net703),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00388_));
 sky130_fd_sc_hd__and2_1 _09758_ (.A(net868),
    .B(net703),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00389_));
 sky130_fd_sc_hd__and2_1 _09759_ (.A(net852),
    .B(net687),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00390_));
 sky130_fd_sc_hd__and2_1 _09760_ (.A(net852),
    .B(net687),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00391_));
 sky130_fd_sc_hd__and2_1 _09761_ (.A(net853),
    .B(net688),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00392_));
 sky130_fd_sc_hd__and2_1 _09762_ (.A(net853),
    .B(net688),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00393_));
 sky130_fd_sc_hd__and2_1 _09763_ (.A(net853),
    .B(net688),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00394_));
 sky130_fd_sc_hd__and2_1 _09764_ (.A(net849),
    .B(net684),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00395_));
 sky130_fd_sc_hd__and2_1 _09765_ (.A(net848),
    .B(net683),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00396_));
 sky130_fd_sc_hd__and2_1 _09766_ (.A(net848),
    .B(net683),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00397_));
 sky130_fd_sc_hd__and2_1 _09767_ (.A(net792),
    .B(net627),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00398_));
 sky130_fd_sc_hd__and2_1 _09768_ (.A(net793),
    .B(net628),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00399_));
 sky130_fd_sc_hd__and2_1 _09769_ (.A(net793),
    .B(net628),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00400_));
 sky130_fd_sc_hd__and2_1 _09770_ (.A(net791),
    .B(net626),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00401_));
 sky130_fd_sc_hd__and2_1 _09771_ (.A(net788),
    .B(net623),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00402_));
 sky130_fd_sc_hd__and2_1 _09772_ (.A(net784),
    .B(net619),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00403_));
 sky130_fd_sc_hd__and2_1 _09773_ (.A(net838),
    .B(net673),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00404_));
 sky130_fd_sc_hd__and2_1 _09774_ (.A(net842),
    .B(net677),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00405_));
 sky130_fd_sc_hd__and2_1 _09775_ (.A(net843),
    .B(net678),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00406_));
 sky130_fd_sc_hd__and2_1 _09776_ (.A(net857),
    .B(net692),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00407_));
 sky130_fd_sc_hd__and2_1 _09777_ (.A(net857),
    .B(net692),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00408_));
 sky130_fd_sc_hd__and2_1 _09778_ (.A(net857),
    .B(net692),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00409_));
 sky130_fd_sc_hd__and2_1 _09779_ (.A(net864),
    .B(net699),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00410_));
 sky130_fd_sc_hd__and2_1 _09780_ (.A(net862),
    .B(net697),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00411_));
 sky130_fd_sc_hd__and2_1 _09781_ (.A(net863),
    .B(net698),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00412_));
 sky130_fd_sc_hd__and2_1 _09782_ (.A(net872),
    .B(net707),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00413_));
 sky130_fd_sc_hd__and2_1 _09783_ (.A(net870),
    .B(net705),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00414_));
 sky130_fd_sc_hd__and2_1 _09784_ (.A(net871),
    .B(net706),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00415_));
 sky130_fd_sc_hd__and2_1 _09785_ (.A(net873),
    .B(net708),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00416_));
 sky130_fd_sc_hd__and2_1 _09786_ (.A(net872),
    .B(net707),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00417_));
 sky130_fd_sc_hd__and2_1 _09787_ (.A(net869),
    .B(net704),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00418_));
 sky130_fd_sc_hd__and2_1 _09788_ (.A(net866),
    .B(net701),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00419_));
 sky130_fd_sc_hd__and2_1 _09789_ (.A(net868),
    .B(net703),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00420_));
 sky130_fd_sc_hd__and2_1 _09790_ (.A(net866),
    .B(net701),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00421_));
 sky130_fd_sc_hd__and2_1 _09791_ (.A(net851),
    .B(net686),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00422_));
 sky130_fd_sc_hd__and2_1 _09792_ (.A(net851),
    .B(net686),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00423_));
 sky130_fd_sc_hd__and2_1 _09793_ (.A(net850),
    .B(net685),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00424_));
 sky130_fd_sc_hd__and2_1 _09794_ (.A(net850),
    .B(net685),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00425_));
 sky130_fd_sc_hd__and2_1 _09795_ (.A(net850),
    .B(net685),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00426_));
 sky130_fd_sc_hd__and2_1 _09796_ (.A(net847),
    .B(net682),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00427_));
 sky130_fd_sc_hd__and2_1 _09797_ (.A(net846),
    .B(net681),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00428_));
 sky130_fd_sc_hd__and2_1 _09798_ (.A(net790),
    .B(net625),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00429_));
 sky130_fd_sc_hd__and2_1 _09799_ (.A(net790),
    .B(net625),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00430_));
 sky130_fd_sc_hd__and2_1 _09800_ (.A(net793),
    .B(net628),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00431_));
 sky130_fd_sc_hd__and2_1 _09801_ (.A(net791),
    .B(net626),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00432_));
 sky130_fd_sc_hd__and2_1 _09802_ (.A(net791),
    .B(net626),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00433_));
 sky130_fd_sc_hd__and2_1 _09803_ (.A(net787),
    .B(net622),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00434_));
 sky130_fd_sc_hd__and2_1 _09804_ (.A(net787),
    .B(net622),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00435_));
 sky130_fd_sc_hd__and2_1 _09805_ (.A(net761),
    .B(net596),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00436_));
 sky130_fd_sc_hd__and2_1 _09806_ (.A(net764),
    .B(net599),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00437_));
 sky130_fd_sc_hd__and2_1 _09807_ (.A(net764),
    .B(net599),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00438_));
 sky130_fd_sc_hd__and2_1 _09808_ (.A(net764),
    .B(net599),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00439_));
 sky130_fd_sc_hd__and2_1 _09809_ (.A(net764),
    .B(net599),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00440_));
 sky130_fd_sc_hd__and2_1 _09810_ (.A(net764),
    .B(net599),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00441_));
 sky130_fd_sc_hd__and2_1 _09811_ (.A(net764),
    .B(net599),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00442_));
 sky130_fd_sc_hd__and2_1 _09812_ (.A(net764),
    .B(net599),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00443_));
 sky130_fd_sc_hd__and2_1 _09813_ (.A(net775),
    .B(net610),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00444_));
 sky130_fd_sc_hd__and2_1 _09814_ (.A(net787),
    .B(net622),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00445_));
 sky130_fd_sc_hd__and2_1 _09815_ (.A(net851),
    .B(net686),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00446_));
 sky130_fd_sc_hd__and2_1 _09816_ (.A(net843),
    .B(net678),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00447_));
 sky130_fd_sc_hd__and2_1 _09817_ (.A(net843),
    .B(net678),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00448_));
 sky130_fd_sc_hd__and2_1 _09818_ (.A(net843),
    .B(net678),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00449_));
 sky130_fd_sc_hd__and2_1 _09819_ (.A(net843),
    .B(net678),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00450_));
 sky130_fd_sc_hd__and2_1 _09820_ (.A(net866),
    .B(net701),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00451_));
 sky130_fd_sc_hd__and2_1 _09821_ (.A(net870),
    .B(net705),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00452_));
 sky130_fd_sc_hd__and2_1 _09822_ (.A(net870),
    .B(net705),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00453_));
 sky130_fd_sc_hd__and2_1 _09823_ (.A(net873),
    .B(net708),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00454_));
 sky130_fd_sc_hd__and2_1 _09824_ (.A(net873),
    .B(net708),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00455_));
 sky130_fd_sc_hd__and2_1 _09825_ (.A(net873),
    .B(net708),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00456_));
 sky130_fd_sc_hd__and2_1 _09826_ (.A(net874),
    .B(net709),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00457_));
 sky130_fd_sc_hd__and2_1 _09827_ (.A(net874),
    .B(net709),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00458_));
 sky130_fd_sc_hd__and2_1 _09828_ (.A(net869),
    .B(net704),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00459_));
 sky130_fd_sc_hd__and2_1 _09829_ (.A(net869),
    .B(net704),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00460_));
 sky130_fd_sc_hd__and2_1 _09830_ (.A(net868),
    .B(net703),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00461_));
 sky130_fd_sc_hd__and2_1 _09831_ (.A(net852),
    .B(net687),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00462_));
 sky130_fd_sc_hd__and2_1 _09832_ (.A(net853),
    .B(net688),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00463_));
 sky130_fd_sc_hd__and2_1 _09833_ (.A(net853),
    .B(net688),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00464_));
 sky130_fd_sc_hd__and2_1 _09834_ (.A(net849),
    .B(net684),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00465_));
 sky130_fd_sc_hd__and2_1 _09835_ (.A(net849),
    .B(net684),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00466_));
 sky130_fd_sc_hd__and2_1 _09836_ (.A(net849),
    .B(net684),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00467_));
 sky130_fd_sc_hd__and2_1 _09837_ (.A(net849),
    .B(net684),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00468_));
 sky130_fd_sc_hd__and2_1 _09838_ (.A(net848),
    .B(net683),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00469_));
 sky130_fd_sc_hd__and2_1 _09839_ (.A(net848),
    .B(net683),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00470_));
 sky130_fd_sc_hd__and2_1 _09840_ (.A(net792),
    .B(net627),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00471_));
 sky130_fd_sc_hd__and2_1 _09841_ (.A(net792),
    .B(net627),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00472_));
 sky130_fd_sc_hd__and2_1 _09842_ (.A(net792),
    .B(net627),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00473_));
 sky130_fd_sc_hd__and2_1 _09843_ (.A(net792),
    .B(net627),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00474_));
 sky130_fd_sc_hd__and2_1 _09844_ (.A(net792),
    .B(net627),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00475_));
 sky130_fd_sc_hd__and2_1 _09845_ (.A(net785),
    .B(net620),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00476_));
 sky130_fd_sc_hd__and2_1 _09846_ (.A(net839),
    .B(net674),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00477_));
 sky130_fd_sc_hd__and2_1 _09847_ (.A(net856),
    .B(net691),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00478_));
 sky130_fd_sc_hd__and2_1 _09848_ (.A(net857),
    .B(net692),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00479_));
 sky130_fd_sc_hd__and2_1 _09849_ (.A(net857),
    .B(net692),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00480_));
 sky130_fd_sc_hd__and2_1 _09850_ (.A(net857),
    .B(net692),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00481_));
 sky130_fd_sc_hd__and2_1 _09851_ (.A(net864),
    .B(net699),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00482_));
 sky130_fd_sc_hd__and2_1 _09852_ (.A(net863),
    .B(net698),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00483_));
 sky130_fd_sc_hd__and2_1 _09853_ (.A(net867),
    .B(net702),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00484_));
 sky130_fd_sc_hd__and2_1 _09854_ (.A(net867),
    .B(net702),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00485_));
 sky130_fd_sc_hd__and2_1 _09855_ (.A(net872),
    .B(net707),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00486_));
 sky130_fd_sc_hd__and2_1 _09856_ (.A(net871),
    .B(net706),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00487_));
 sky130_fd_sc_hd__and2_1 _09857_ (.A(net871),
    .B(net706),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00488_));
 sky130_fd_sc_hd__and2_1 _09858_ (.A(net872),
    .B(net707),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00489_));
 sky130_fd_sc_hd__and2_1 _09859_ (.A(net867),
    .B(net702),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00490_));
 sky130_fd_sc_hd__and2_1 _09860_ (.A(net866),
    .B(net701),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00491_));
 sky130_fd_sc_hd__and2_1 _09861_ (.A(net867),
    .B(net702),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00492_));
 sky130_fd_sc_hd__and2_1 _09862_ (.A(net866),
    .B(net701),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00493_));
 sky130_fd_sc_hd__and2_1 _09863_ (.A(net851),
    .B(net686),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00494_));
 sky130_fd_sc_hd__and2_1 _09864_ (.A(net851),
    .B(net686),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00495_));
 sky130_fd_sc_hd__and2_1 _09865_ (.A(net850),
    .B(net685),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00496_));
 sky130_fd_sc_hd__and2_1 _09866_ (.A(net850),
    .B(net685),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00497_));
 sky130_fd_sc_hd__and2_1 _09867_ (.A(net847),
    .B(net682),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00498_));
 sky130_fd_sc_hd__and2_1 _09868_ (.A(net847),
    .B(net682),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00499_));
 sky130_fd_sc_hd__and2_1 _09869_ (.A(net847),
    .B(net682),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00500_));
 sky130_fd_sc_hd__and2_1 _09870_ (.A(net846),
    .B(net681),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00501_));
 sky130_fd_sc_hd__and2_1 _09871_ (.A(net846),
    .B(net681),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00502_));
 sky130_fd_sc_hd__and2_1 _09872_ (.A(net790),
    .B(net625),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00503_));
 sky130_fd_sc_hd__and2_1 _09873_ (.A(net790),
    .B(net625),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00504_));
 sky130_fd_sc_hd__and2_1 _09874_ (.A(net790),
    .B(net625),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00505_));
 sky130_fd_sc_hd__and2_1 _09875_ (.A(net791),
    .B(net626),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00506_));
 sky130_fd_sc_hd__and2_1 _09876_ (.A(net846),
    .B(net681),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00507_));
 sky130_fd_sc_hd__and2_1 _09877_ (.A(net846),
    .B(net681),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00508_));
 sky130_fd_sc_hd__and2_1 _09878_ (.A(net847),
    .B(net682),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00509_));
 sky130_fd_sc_hd__and2_1 _09879_ (.A(net866),
    .B(net701),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00510_));
 sky130_fd_sc_hd__and2_1 _09880_ (.A(net858),
    .B(net693),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00511_));
 sky130_fd_sc_hd__and2_1 _09881_ (.A(net858),
    .B(net693),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00512_));
 sky130_fd_sc_hd__and2_1 _09882_ (.A(net856),
    .B(net691),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00513_));
 sky130_fd_sc_hd__and2_1 _09883_ (.A(net866),
    .B(net701),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00514_));
 sky130_fd_sc_hd__and2_1 _09884_ (.A(net867),
    .B(net702),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00515_));
 sky130_fd_sc_hd__and2_1 _09885_ (.A(net870),
    .B(net705),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00516_));
 sky130_fd_sc_hd__and2_1 _09886_ (.A(net872),
    .B(net707),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00517_));
 sky130_fd_sc_hd__and2_1 _09887_ (.A(net873),
    .B(net708),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00518_));
 sky130_fd_sc_hd__and2_1 _09888_ (.A(net875),
    .B(net710),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00519_));
 sky130_fd_sc_hd__and2_1 _09889_ (.A(net875),
    .B(net710),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00520_));
 sky130_fd_sc_hd__and2_1 _09890_ (.A(net874),
    .B(net709),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00521_));
 sky130_fd_sc_hd__and2_1 _09891_ (.A(net874),
    .B(net709),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00522_));
 sky130_fd_sc_hd__and2_1 _09892_ (.A(net874),
    .B(net709),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00523_));
 sky130_fd_sc_hd__and2_1 _09893_ (.A(net869),
    .B(net704),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00524_));
 sky130_fd_sc_hd__and2_1 _09894_ (.A(net868),
    .B(net703),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00525_));
 sky130_fd_sc_hd__and2_1 _09895_ (.A(net868),
    .B(net703),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00526_));
 sky130_fd_sc_hd__and2_1 _09896_ (.A(net852),
    .B(net687),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00527_));
 sky130_fd_sc_hd__and2_1 _09897_ (.A(net852),
    .B(net687),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00528_));
 sky130_fd_sc_hd__and2_1 _09898_ (.A(net854),
    .B(net689),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00529_));
 sky130_fd_sc_hd__and2_1 _09899_ (.A(net853),
    .B(net688),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00530_));
 sky130_fd_sc_hd__and2_1 _09900_ (.A(net853),
    .B(net688),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00531_));
 sky130_fd_sc_hd__and2_1 _09901_ (.A(net848),
    .B(net683),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00532_));
 sky130_fd_sc_hd__and2_1 _09902_ (.A(net793),
    .B(net628),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00533_));
 sky130_fd_sc_hd__and2_1 _09903_ (.A(net793),
    .B(net628),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00534_));
 sky130_fd_sc_hd__and2_1 _09904_ (.A(net793),
    .B(net628),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00535_));
 sky130_fd_sc_hd__and2_1 _09905_ (.A(net789),
    .B(net624),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00536_));
 sky130_fd_sc_hd__and2_1 _09906_ (.A(net793),
    .B(net628),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00537_));
 sky130_fd_sc_hd__and2_1 _09907_ (.A(net793),
    .B(net628),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00538_));
 sky130_fd_sc_hd__and2_1 _09908_ (.A(net789),
    .B(net624),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00539_));
 sky130_fd_sc_hd__and2_1 _09909_ (.A(net784),
    .B(net619),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00540_));
 sky130_fd_sc_hd__and2_1 _09910_ (.A(net839),
    .B(net674),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00541_));
 sky130_fd_sc_hd__and2_1 _09911_ (.A(net864),
    .B(net699),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00542_));
 sky130_fd_sc_hd__and2_1 _09912_ (.A(net857),
    .B(net692),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00543_));
 sky130_fd_sc_hd__and2_1 _09913_ (.A(net858),
    .B(net693),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00544_));
 sky130_fd_sc_hd__and2_1 _09914_ (.A(net864),
    .B(net699),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00545_));
 sky130_fd_sc_hd__and2_1 _09915_ (.A(net864),
    .B(net699),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00546_));
 sky130_fd_sc_hd__and2_1 _09916_ (.A(net864),
    .B(net699),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00547_));
 sky130_fd_sc_hd__and2_1 _09917_ (.A(net864),
    .B(net699),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00548_));
 sky130_fd_sc_hd__and2_1 _09918_ (.A(net872),
    .B(net707),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00549_));
 sky130_fd_sc_hd__and2_1 _09919_ (.A(net871),
    .B(net706),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00550_));
 sky130_fd_sc_hd__and2_1 _09920_ (.A(net871),
    .B(net706),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00551_));
 sky130_fd_sc_hd__and2_1 _09921_ (.A(net873),
    .B(net708),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00552_));
 sky130_fd_sc_hd__and2_1 _09922_ (.A(net874),
    .B(net709),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00553_));
 sky130_fd_sc_hd__and2_1 _09923_ (.A(net874),
    .B(net709),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00554_));
 sky130_fd_sc_hd__and2_1 _09924_ (.A(net869),
    .B(net704),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00555_));
 sky130_fd_sc_hd__and2_1 _09925_ (.A(net868),
    .B(net703),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00556_));
 sky130_fd_sc_hd__and2_1 _09926_ (.A(net852),
    .B(net687),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00557_));
 sky130_fd_sc_hd__and2_1 _09927_ (.A(net852),
    .B(net687),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00558_));
 sky130_fd_sc_hd__and2_1 _09928_ (.A(net852),
    .B(net687),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00559_));
 sky130_fd_sc_hd__and2_1 _09929_ (.A(net850),
    .B(net685),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00560_));
 sky130_fd_sc_hd__and2_1 _09930_ (.A(net850),
    .B(net685),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00561_));
 sky130_fd_sc_hd__and2_1 _09931_ (.A(net847),
    .B(net682),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00562_));
 sky130_fd_sc_hd__and2_1 _09932_ (.A(net847),
    .B(net682),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00563_));
 sky130_fd_sc_hd__and2_1 _09933_ (.A(net846),
    .B(net681),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00564_));
 sky130_fd_sc_hd__and2_1 _09934_ (.A(net790),
    .B(net625),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00565_));
 sky130_fd_sc_hd__and2_1 _09935_ (.A(net794),
    .B(net629),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00566_));
 sky130_fd_sc_hd__and2_1 _09936_ (.A(net793),
    .B(net628),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00567_));
 sky130_fd_sc_hd__and2_1 _09937_ (.A(net791),
    .B(net626),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00568_));
 sky130_fd_sc_hd__and2_1 _09938_ (.A(net791),
    .B(net626),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00569_));
 sky130_fd_sc_hd__and2_1 _09939_ (.A(net791),
    .B(net626),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00570_));
 sky130_fd_sc_hd__and2_1 _09940_ (.A(net788),
    .B(net623),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00571_));
 sky130_fd_sc_hd__and2_1 _09941_ (.A(net788),
    .B(net623),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00572_));
 sky130_fd_sc_hd__and2_1 _09942_ (.A(net794),
    .B(net629),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00573_));
 sky130_fd_sc_hd__and2_1 _09943_ (.A(net789),
    .B(net624),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00574_));
 sky130_fd_sc_hd__and2_1 _09944_ (.A(net789),
    .B(net624),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00575_));
 sky130_fd_sc_hd__and2_1 _09945_ (.A(net789),
    .B(net624),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00576_));
 sky130_fd_sc_hd__and2_1 _09946_ (.A(net789),
    .B(net624),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00577_));
 sky130_fd_sc_hd__and2_1 _09947_ (.A(net794),
    .B(net629),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00578_));
 sky130_fd_sc_hd__and2_1 _09948_ (.A(net789),
    .B(net624),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00579_));
 sky130_fd_sc_hd__and2_1 _09949_ (.A(net767),
    .B(net602),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00580_));
 sky130_fd_sc_hd__and2_1 _09950_ (.A(net768),
    .B(net603),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00581_));
 sky130_fd_sc_hd__and2_1 _09951_ (.A(net767),
    .B(net602),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00582_));
 sky130_fd_sc_hd__and2_1 _09952_ (.A(net767),
    .B(net602),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00583_));
 sky130_fd_sc_hd__and2_1 _09953_ (.A(net771),
    .B(net606),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00584_));
 sky130_fd_sc_hd__and2_1 _09954_ (.A(net771),
    .B(net606),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00585_));
 sky130_fd_sc_hd__and2_1 _09955_ (.A(net771),
    .B(net606),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00586_));
 sky130_fd_sc_hd__and2_1 _09956_ (.A(net772),
    .B(net607),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00587_));
 sky130_fd_sc_hd__and2_1 _09957_ (.A(net773),
    .B(net608),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00588_));
 sky130_fd_sc_hd__and2_1 _09958_ (.A(net770),
    .B(net605),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00589_));
 sky130_fd_sc_hd__and2_1 _09959_ (.A(net775),
    .B(net610),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00590_));
 sky130_fd_sc_hd__and2_1 _09960_ (.A(net770),
    .B(net605),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00591_));
 sky130_fd_sc_hd__and2_1 _09961_ (.A(net775),
    .B(net610),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00592_));
 sky130_fd_sc_hd__and2_1 _09962_ (.A(net775),
    .B(net610),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00593_));
 sky130_fd_sc_hd__and2_1 _09963_ (.A(net775),
    .B(net610),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00594_));
 sky130_fd_sc_hd__and2_1 _09964_ (.A(net775),
    .B(net610),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00595_));
 sky130_fd_sc_hd__and2_1 _09965_ (.A(net773),
    .B(net608),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00596_));
 sky130_fd_sc_hd__and2_1 _09966_ (.A(net772),
    .B(net607),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00597_));
 sky130_fd_sc_hd__and2_1 _09967_ (.A(net773),
    .B(net608),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00598_));
 sky130_fd_sc_hd__and2_1 _09968_ (.A(net751),
    .B(net586),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00599_));
 sky130_fd_sc_hd__and2_1 _09969_ (.A(net751),
    .B(net586),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00600_));
 sky130_fd_sc_hd__and2_1 _09970_ (.A(net751),
    .B(net586),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00601_));
 sky130_fd_sc_hd__and2_1 _09971_ (.A(net750),
    .B(net585),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00602_));
 sky130_fd_sc_hd__and2_1 _09972_ (.A(net754),
    .B(net589),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00603_));
 sky130_fd_sc_hd__and2_1 _09973_ (.A(net782),
    .B(net617),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00604_));
 sky130_fd_sc_hd__and2_1 _09974_ (.A(net782),
    .B(net617),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00605_));
 sky130_fd_sc_hd__and2_1 _09975_ (.A(net782),
    .B(net617),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00606_));
 sky130_fd_sc_hd__and2_1 _09976_ (.A(net782),
    .B(net617),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00607_));
 sky130_fd_sc_hd__and2_1 _09977_ (.A(net782),
    .B(net617),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00608_));
 sky130_fd_sc_hd__and2_1 _09978_ (.A(net782),
    .B(net617),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00609_));
 sky130_fd_sc_hd__and2_1 _09979_ (.A(net783),
    .B(net618),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00610_));
 sky130_fd_sc_hd__and2_1 _09980_ (.A(net754),
    .B(net589),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00611_));
 sky130_fd_sc_hd__and2_1 _09981_ (.A(net755),
    .B(net590),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00612_));
 sky130_fd_sc_hd__and2_1 _09982_ (.A(net751),
    .B(net586),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00613_));
 sky130_fd_sc_hd__and2_1 _09983_ (.A(net832),
    .B(net667),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00614_));
 sky130_fd_sc_hd__and2_1 _09984_ (.A(net831),
    .B(net666),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00615_));
 sky130_fd_sc_hd__and2_1 _09985_ (.A(net831),
    .B(net666),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00616_));
 sky130_fd_sc_hd__and2_1 _09986_ (.A(net831),
    .B(net666),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00617_));
 sky130_fd_sc_hd__and2_1 _09987_ (.A(net831),
    .B(net666),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00618_));
 sky130_fd_sc_hd__and2_1 _09988_ (.A(net831),
    .B(net666),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00619_));
 sky130_fd_sc_hd__and2_1 _09989_ (.A(net832),
    .B(net667),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00620_));
 sky130_fd_sc_hd__and2_1 _09990_ (.A(net831),
    .B(net666),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00621_));
 sky130_fd_sc_hd__and2_1 _09991_ (.A(net860),
    .B(net695),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00622_));
 sky130_fd_sc_hd__and2_1 _09992_ (.A(net832),
    .B(net667),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00623_));
 sky130_fd_sc_hd__and2_1 _09993_ (.A(net832),
    .B(net667),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00624_));
 sky130_fd_sc_hd__and2_1 _09994_ (.A(net860),
    .B(net695),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00625_));
 sky130_fd_sc_hd__and2_1 _09995_ (.A(net860),
    .B(net695),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00626_));
 sky130_fd_sc_hd__and2_1 _09996_ (.A(net861),
    .B(net696),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00627_));
 sky130_fd_sc_hd__and2_1 _09997_ (.A(net861),
    .B(net696),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00628_));
 sky130_fd_sc_hd__and2_1 _09998_ (.A(net861),
    .B(net696),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00629_));
 sky130_fd_sc_hd__and2_1 _09999_ (.A(net855),
    .B(net690),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00630_));
 sky130_fd_sc_hd__and2_1 _10000_ (.A(net855),
    .B(net690),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00631_));
 sky130_fd_sc_hd__and2_1 _10001_ (.A(net855),
    .B(net690),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00632_));
 sky130_fd_sc_hd__and2_1 _10002_ (.A(net813),
    .B(net648),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00633_));
 sky130_fd_sc_hd__and2_1 _10003_ (.A(net814),
    .B(net649),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00634_));
 sky130_fd_sc_hd__and2_1 _10004_ (.A(net840),
    .B(net675),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00635_));
 sky130_fd_sc_hd__and2_1 _10005_ (.A(net841),
    .B(net676),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00636_));
 sky130_fd_sc_hd__and2_1 _10006_ (.A(net814),
    .B(net649),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00637_));
 sky130_fd_sc_hd__and2_1 _10007_ (.A(net813),
    .B(net648),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00638_));
 sky130_fd_sc_hd__and2_1 _10008_ (.A(net840),
    .B(net675),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00639_));
 sky130_fd_sc_hd__and2_1 _10009_ (.A(net811),
    .B(net646),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00640_));
 sky130_fd_sc_hd__and2_1 _10010_ (.A(net811),
    .B(net646),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00641_));
 sky130_fd_sc_hd__and2_1 _10011_ (.A(net811),
    .B(net646),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00642_));
 sky130_fd_sc_hd__and2_1 _10012_ (.A(net809),
    .B(net644),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00643_));
 sky130_fd_sc_hd__and2_1 _10013_ (.A(net811),
    .B(net646),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00644_));
 sky130_fd_sc_hd__and2_1 _10014_ (.A(net809),
    .B(net644),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00645_));
 sky130_fd_sc_hd__and2_1 _10015_ (.A(net827),
    .B(net662),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00646_));
 sky130_fd_sc_hd__and2_1 _10016_ (.A(net830),
    .B(net665),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00647_));
 sky130_fd_sc_hd__and2_1 _10017_ (.A(net827),
    .B(net662),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00648_));
 sky130_fd_sc_hd__and2_1 _10018_ (.A(net827),
    .B(net662),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00649_));
 sky130_fd_sc_hd__and2_1 _10019_ (.A(net827),
    .B(net662),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00650_));
 sky130_fd_sc_hd__and2_1 _10020_ (.A(net830),
    .B(net665),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00651_));
 sky130_fd_sc_hd__and2_1 _10021_ (.A(net830),
    .B(net665),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00652_));
 sky130_fd_sc_hd__and2_1 _10022_ (.A(net830),
    .B(net665),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00653_));
 sky130_fd_sc_hd__and2_1 _10023_ (.A(net855),
    .B(net690),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00654_));
 sky130_fd_sc_hd__and2_1 _10024_ (.A(net829),
    .B(net664),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00655_));
 sky130_fd_sc_hd__and2_1 _10025_ (.A(net833),
    .B(net668),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00656_));
 sky130_fd_sc_hd__and2_1 _10026_ (.A(net859),
    .B(net694),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00657_));
 sky130_fd_sc_hd__and2_1 _10027_ (.A(net855),
    .B(net690),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00658_));
 sky130_fd_sc_hd__and2_1 _10028_ (.A(net855),
    .B(net690),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00659_));
 sky130_fd_sc_hd__and2_1 _10029_ (.A(net839),
    .B(net674),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00660_));
 sky130_fd_sc_hd__and2_1 _10030_ (.A(net785),
    .B(net620),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00661_));
 sky130_fd_sc_hd__and2_1 _10031_ (.A(net783),
    .B(net618),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00662_));
 sky130_fd_sc_hd__and2_1 _10032_ (.A(net836),
    .B(net671),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00663_));
 sky130_fd_sc_hd__and2_1 _10033_ (.A(net836),
    .B(net671),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00664_));
 sky130_fd_sc_hd__and2_1 _10034_ (.A(net785),
    .B(net620),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00665_));
 sky130_fd_sc_hd__and2_1 _10035_ (.A(net836),
    .B(net671),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00666_));
 sky130_fd_sc_hd__and2_1 _10036_ (.A(net836),
    .B(net671),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00667_));
 sky130_fd_sc_hd__and2_1 _10037_ (.A(net756),
    .B(net591),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00668_));
 sky130_fd_sc_hd__and2_1 _10038_ (.A(net837),
    .B(net672),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00669_));
 sky130_fd_sc_hd__and2_1 _10039_ (.A(net838),
    .B(net673),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00670_));
 sky130_fd_sc_hd__and2_1 _10040_ (.A(net836),
    .B(net671),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00671_));
 sky130_fd_sc_hd__and2_1 _10041_ (.A(net836),
    .B(net671),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00672_));
 sky130_fd_sc_hd__and2_1 _10042_ (.A(net836),
    .B(net671),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00673_));
 sky130_fd_sc_hd__and2_1 _10043_ (.A(net838),
    .B(net673),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00674_));
 sky130_fd_sc_hd__and2_1 _10044_ (.A(net783),
    .B(net618),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00675_));
 sky130_fd_sc_hd__and2_1 _10045_ (.A(net782),
    .B(net617),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00676_));
 sky130_fd_sc_hd__and2_1 _10046_ (.A(net811),
    .B(net646),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00677_));
 sky130_fd_sc_hd__and2_1 _10047_ (.A(net756),
    .B(net591),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00678_));
 sky130_fd_sc_hd__and2_1 _10048_ (.A(net761),
    .B(net596),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00679_));
 sky130_fd_sc_hd__and2_1 _10049_ (.A(net759),
    .B(net594),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00680_));
 sky130_fd_sc_hd__and2_1 _10050_ (.A(net761),
    .B(net596),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00681_));
 sky130_fd_sc_hd__and2_1 _10051_ (.A(net764),
    .B(net599),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00682_));
 sky130_fd_sc_hd__and2_1 _10052_ (.A(net764),
    .B(net599),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00683_));
 sky130_fd_sc_hd__and2_1 _10053_ (.A(net759),
    .B(net594),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00684_));
 sky130_fd_sc_hd__and2_1 _10054_ (.A(net761),
    .B(net596),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00685_));
 sky130_fd_sc_hd__and2_1 _10055_ (.A(net719),
    .B(net554),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00686_));
 sky130_fd_sc_hd__and2_1 _10056_ (.A(net719),
    .B(net554),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00687_));
 sky130_fd_sc_hd__and2_1 _10057_ (.A(net719),
    .B(net554),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00688_));
 sky130_fd_sc_hd__and2_1 _10058_ (.A(net719),
    .B(net554),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00689_));
 sky130_fd_sc_hd__and2_1 _10059_ (.A(net719),
    .B(net554),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00690_));
 sky130_fd_sc_hd__and2_1 _10060_ (.A(net720),
    .B(net555),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00691_));
 sky130_fd_sc_hd__and2_1 _10061_ (.A(net720),
    .B(net555),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00692_));
 sky130_fd_sc_hd__and2_1 _10062_ (.A(net720),
    .B(net555),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00693_));
 sky130_fd_sc_hd__and2_1 _10063_ (.A(net783),
    .B(net618),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00694_));
 sky130_fd_sc_hd__and2_1 _10064_ (.A(net783),
    .B(net618),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00695_));
 sky130_fd_sc_hd__and2_1 _10065_ (.A(net783),
    .B(net618),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00696_));
 sky130_fd_sc_hd__and2_1 _10066_ (.A(net783),
    .B(net618),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00697_));
 sky130_fd_sc_hd__and2_1 _10067_ (.A(net783),
    .B(net618),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00698_));
 sky130_fd_sc_hd__and2_1 _10068_ (.A(net782),
    .B(net617),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00699_));
 sky130_fd_sc_hd__and2_1 _10069_ (.A(net783),
    .B(net618),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00700_));
 sky130_fd_sc_hd__and2_1 _10070_ (.A(net756),
    .B(net591),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00701_));
 sky130_fd_sc_hd__and2_1 _10071_ (.A(net756),
    .B(net591),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00702_));
 sky130_fd_sc_hd__and2_1 _10072_ (.A(net784),
    .B(net619),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00703_));
 sky130_fd_sc_hd__and2_1 _10073_ (.A(net784),
    .B(net619),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00704_));
 sky130_fd_sc_hd__and2_1 _10074_ (.A(net786),
    .B(net621),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00705_));
 sky130_fd_sc_hd__and2_1 _10075_ (.A(net836),
    .B(net671),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00706_));
 sky130_fd_sc_hd__and2_1 _10076_ (.A(net836),
    .B(net671),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00707_));
 sky130_fd_sc_hd__and2_1 _10077_ (.A(net784),
    .B(net619),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00708_));
 sky130_fd_sc_hd__and2_1 _10078_ (.A(net786),
    .B(net621),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00709_));
 sky130_fd_sc_hd__and2_1 _10079_ (.A(net756),
    .B(net591),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00710_));
 sky130_fd_sc_hd__and2_1 _10080_ (.A(net757),
    .B(net592),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00711_));
 sky130_fd_sc_hd__and2_1 _10081_ (.A(net822),
    .B(net657),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00712_));
 sky130_fd_sc_hd__and2_1 _10082_ (.A(net822),
    .B(net657),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00713_));
 sky130_fd_sc_hd__and2_1 _10083_ (.A(net822),
    .B(net657),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00714_));
 sky130_fd_sc_hd__and2_1 _10084_ (.A(net822),
    .B(net657),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00715_));
 sky130_fd_sc_hd__and2_1 _10085_ (.A(net822),
    .B(net657),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00716_));
 sky130_fd_sc_hd__and2_1 _10086_ (.A(net823),
    .B(net658),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00717_));
 sky130_fd_sc_hd__and2_1 _10087_ (.A(net823),
    .B(net658),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00718_));
 sky130_fd_sc_hd__and2_1 _10088_ (.A(net824),
    .B(net659),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00719_));
 sky130_fd_sc_hd__and2_1 _10089_ (.A(net832),
    .B(net667),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00720_));
 sky130_fd_sc_hd__and2_1 _10090_ (.A(net831),
    .B(net666),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00721_));
 sky130_fd_sc_hd__and2_1 _10091_ (.A(net834),
    .B(net669),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00722_));
 sky130_fd_sc_hd__and2_1 _10092_ (.A(net831),
    .B(net666),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00723_));
 sky130_fd_sc_hd__and2_1 _10093_ (.A(net833),
    .B(net668),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00724_));
 sky130_fd_sc_hd__and2_1 _10094_ (.A(net831),
    .B(net666),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00725_));
 sky130_fd_sc_hd__and2_1 _10095_ (.A(net833),
    .B(net668),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00726_));
 sky130_fd_sc_hd__and2_1 _10096_ (.A(net827),
    .B(net662),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00727_));
 sky130_fd_sc_hd__and2_1 _10097_ (.A(net814),
    .B(net649),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00728_));
 sky130_fd_sc_hd__and2_1 _10098_ (.A(net830),
    .B(net665),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00729_));
 sky130_fd_sc_hd__and2_1 _10099_ (.A(net814),
    .B(net649),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00730_));
 sky130_fd_sc_hd__and2_1 _10100_ (.A(net814),
    .B(net649),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00731_));
 sky130_fd_sc_hd__and2_1 _10101_ (.A(net814),
    .B(net649),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00732_));
 sky130_fd_sc_hd__and2_1 _10102_ (.A(net814),
    .B(net649),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00733_));
 sky130_fd_sc_hd__and2_1 _10103_ (.A(net814),
    .B(net649),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00734_));
 sky130_fd_sc_hd__and2_1 _10104_ (.A(net813),
    .B(net648),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00735_));
 sky130_fd_sc_hd__and2_1 _10105_ (.A(net811),
    .B(net646),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00736_));
 sky130_fd_sc_hd__and2_1 _10106_ (.A(net811),
    .B(net646),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00737_));
 sky130_fd_sc_hd__and2_1 _10107_ (.A(net812),
    .B(net647),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00738_));
 sky130_fd_sc_hd__and2_1 _10108_ (.A(net810),
    .B(net645),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00739_));
 sky130_fd_sc_hd__and2_1 _10109_ (.A(net809),
    .B(net644),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00740_));
 sky130_fd_sc_hd__and2_1 _10110_ (.A(net809),
    .B(net644),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00741_));
 sky130_fd_sc_hd__and2_1 _10111_ (.A(net809),
    .B(net644),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00742_));
 sky130_fd_sc_hd__and2_1 _10112_ (.A(net809),
    .B(net644),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00743_));
 sky130_fd_sc_hd__and2_1 _10113_ (.A(net806),
    .B(net641),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00744_));
 sky130_fd_sc_hd__and2_1 _10114_ (.A(net802),
    .B(net637),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00745_));
 sky130_fd_sc_hd__and2_1 _10115_ (.A(net806),
    .B(net641),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00746_));
 sky130_fd_sc_hd__and2_1 _10116_ (.A(net806),
    .B(net641),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00747_));
 sky130_fd_sc_hd__and2_1 _10117_ (.A(net806),
    .B(net641),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00748_));
 sky130_fd_sc_hd__and2_1 _10118_ (.A(net806),
    .B(net641),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00749_));
 sky130_fd_sc_hd__and2_1 _10119_ (.A(net806),
    .B(net641),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00750_));
 sky130_fd_sc_hd__and2_1 _10120_ (.A(net806),
    .B(net641),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00751_));
 sky130_fd_sc_hd__and2_1 _10121_ (.A(net829),
    .B(net664),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00752_));
 sky130_fd_sc_hd__and2_1 _10122_ (.A(net817),
    .B(net652),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00753_));
 sky130_fd_sc_hd__and2_1 _10123_ (.A(net833),
    .B(net668),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00754_));
 sky130_fd_sc_hd__and2_1 _10124_ (.A(net819),
    .B(net654),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00755_));
 sky130_fd_sc_hd__and2_1 _10125_ (.A(net820),
    .B(net655),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00756_));
 sky130_fd_sc_hd__and2_1 _10126_ (.A(net819),
    .B(net654),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00757_));
 sky130_fd_sc_hd__and2_1 _10127_ (.A(net781),
    .B(net616),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00758_));
 sky130_fd_sc_hd__and2_1 _10128_ (.A(net779),
    .B(net614),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00759_));
 sky130_fd_sc_hd__and2_1 _10129_ (.A(net781),
    .B(net616),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00760_));
 sky130_fd_sc_hd__and2_1 _10130_ (.A(net781),
    .B(net616),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00761_));
 sky130_fd_sc_hd__and2_1 _10131_ (.A(net781),
    .B(net616),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00762_));
 sky130_fd_sc_hd__and2_1 _10132_ (.A(net781),
    .B(net616),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00763_));
 sky130_fd_sc_hd__and2_1 _10133_ (.A(net781),
    .B(net616),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00764_));
 sky130_fd_sc_hd__and2_1 _10134_ (.A(net752),
    .B(net587),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00765_));
 sky130_fd_sc_hd__and2_1 _10135_ (.A(net778),
    .B(net613),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00766_));
 sky130_fd_sc_hd__and2_1 _10136_ (.A(net779),
    .B(net614),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00767_));
 sky130_fd_sc_hd__and2_1 _10137_ (.A(net779),
    .B(net614),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00768_));
 sky130_fd_sc_hd__and2_1 _10138_ (.A(net778),
    .B(net613),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00769_));
 sky130_fd_sc_hd__and2_1 _10139_ (.A(net781),
    .B(net616),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00770_));
 sky130_fd_sc_hd__and2_1 _10140_ (.A(net763),
    .B(net598),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00771_));
 sky130_fd_sc_hd__and2_1 _10141_ (.A(net763),
    .B(net598),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00772_));
 sky130_fd_sc_hd__and2_1 _10142_ (.A(net735),
    .B(net570),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00773_));
 sky130_fd_sc_hd__and2_1 _10143_ (.A(net781),
    .B(net616),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00774_));
 sky130_fd_sc_hd__and2_1 _10144_ (.A(net781),
    .B(net616),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00775_));
 sky130_fd_sc_hd__and2_1 _10145_ (.A(net782),
    .B(net617),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00776_));
 sky130_fd_sc_hd__and2_1 _10146_ (.A(net782),
    .B(net617),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00777_));
 sky130_fd_sc_hd__and2_1 _10147_ (.A(net781),
    .B(net616),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00778_));
 sky130_fd_sc_hd__and2_1 _10148_ (.A(net756),
    .B(net591),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00779_));
 sky130_fd_sc_hd__and2_1 _10149_ (.A(net756),
    .B(net591),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00780_));
 sky130_fd_sc_hd__and2_1 _10150_ (.A(net752),
    .B(net587),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00781_));
 sky130_fd_sc_hd__and2_1 _10151_ (.A(net753),
    .B(net588),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00782_));
 sky130_fd_sc_hd__and2_1 _10152_ (.A(net751),
    .B(net586),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00783_));
 sky130_fd_sc_hd__and2_1 _10153_ (.A(net753),
    .B(net588),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00784_));
 sky130_fd_sc_hd__and2_1 _10154_ (.A(net752),
    .B(net587),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00785_));
 sky130_fd_sc_hd__and2_1 _10155_ (.A(net821),
    .B(net656),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00786_));
 sky130_fd_sc_hd__and2_1 _10156_ (.A(net821),
    .B(net656),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00787_));
 sky130_fd_sc_hd__and2_1 _10157_ (.A(net821),
    .B(net656),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00788_));
 sky130_fd_sc_hd__and2_1 _10158_ (.A(net821),
    .B(net656),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00789_));
 sky130_fd_sc_hd__and2_1 _10159_ (.A(net821),
    .B(net656),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00790_));
 sky130_fd_sc_hd__and2_1 _10160_ (.A(net821),
    .B(net656),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00791_));
 sky130_fd_sc_hd__and2_1 _10161_ (.A(net821),
    .B(net656),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00792_));
 sky130_fd_sc_hd__and2_1 _10162_ (.A(net823),
    .B(net658),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00793_));
 sky130_fd_sc_hd__and2_1 _10163_ (.A(net823),
    .B(net658),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00794_));
 sky130_fd_sc_hd__and2_1 _10164_ (.A(net823),
    .B(net658),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00795_));
 sky130_fd_sc_hd__and2_1 _10165_ (.A(net823),
    .B(net658),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00796_));
 sky130_fd_sc_hd__and2_1 _10166_ (.A(net823),
    .B(net658),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00797_));
 sky130_fd_sc_hd__and2_1 _10167_ (.A(net820),
    .B(net655),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00798_));
 sky130_fd_sc_hd__and2_1 _10168_ (.A(net820),
    .B(net655),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00799_));
 sky130_fd_sc_hd__and2_1 _10169_ (.A(net827),
    .B(net662),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00800_));
 sky130_fd_sc_hd__and2_1 _10170_ (.A(net827),
    .B(net662),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00801_));
 sky130_fd_sc_hd__and2_1 _10171_ (.A(net806),
    .B(net641),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00802_));
 sky130_fd_sc_hd__and2_1 _10172_ (.A(net807),
    .B(net642),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00803_));
 sky130_fd_sc_hd__and2_1 _10173_ (.A(net815),
    .B(net650),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00804_));
 sky130_fd_sc_hd__and2_1 _10174_ (.A(net815),
    .B(net650),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00805_));
 sky130_fd_sc_hd__and2_1 _10175_ (.A(net815),
    .B(net650),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00806_));
 sky130_fd_sc_hd__and2_1 _10176_ (.A(net815),
    .B(net650),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00807_));
 sky130_fd_sc_hd__and2_1 _10177_ (.A(net813),
    .B(net648),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00808_));
 sky130_fd_sc_hd__and2_1 _10178_ (.A(net813),
    .B(net648),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00809_));
 sky130_fd_sc_hd__and2_1 _10179_ (.A(net810),
    .B(net645),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00810_));
 sky130_fd_sc_hd__and2_1 _10180_ (.A(net812),
    .B(net647),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00811_));
 sky130_fd_sc_hd__and2_1 _10181_ (.A(net809),
    .B(net644),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00812_));
 sky130_fd_sc_hd__and2_1 _10182_ (.A(net809),
    .B(net644),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00813_));
 sky130_fd_sc_hd__and2_1 _10183_ (.A(net802),
    .B(net637),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00814_));
 sky130_fd_sc_hd__and2_1 _10184_ (.A(net801),
    .B(net636),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00815_));
 sky130_fd_sc_hd__and2_1 _10185_ (.A(net802),
    .B(net637),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00816_));
 sky130_fd_sc_hd__and2_1 _10186_ (.A(net802),
    .B(net637),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00817_));
 sky130_fd_sc_hd__and2_1 _10187_ (.A(net802),
    .B(net637),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00818_));
 sky130_fd_sc_hd__and2_1 _10188_ (.A(net800),
    .B(net635),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00819_));
 sky130_fd_sc_hd__and2_1 _10189_ (.A(net799),
    .B(net634),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00820_));
 sky130_fd_sc_hd__and2_1 _10190_ (.A(net804),
    .B(net639),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00821_));
 sky130_fd_sc_hd__and2_1 _10191_ (.A(net804),
    .B(net639),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00822_));
 sky130_fd_sc_hd__and2_1 _10192_ (.A(net804),
    .B(net639),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00823_));
 sky130_fd_sc_hd__and2_1 _10193_ (.A(net804),
    .B(net639),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00824_));
 sky130_fd_sc_hd__and2_1 _10194_ (.A(net804),
    .B(net639),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00825_));
 sky130_fd_sc_hd__and2_1 _10195_ (.A(net805),
    .B(net640),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00826_));
 sky130_fd_sc_hd__and2_1 _10196_ (.A(net817),
    .B(net652),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00827_));
 sky130_fd_sc_hd__and2_1 _10197_ (.A(net817),
    .B(net652),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00828_));
 sky130_fd_sc_hd__and2_1 _10198_ (.A(net817),
    .B(net652),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00829_));
 sky130_fd_sc_hd__and2_1 _10199_ (.A(net819),
    .B(net654),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00830_));
 sky130_fd_sc_hd__and2_1 _10200_ (.A(net819),
    .B(net654),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00831_));
 sky130_fd_sc_hd__and2_1 _10201_ (.A(net754),
    .B(net589),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00832_));
 sky130_fd_sc_hd__and2_1 _10202_ (.A(net825),
    .B(net660),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00833_));
 sky130_fd_sc_hd__and2_1 _10203_ (.A(net821),
    .B(net656),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00834_));
 sky130_fd_sc_hd__and2_1 _10204_ (.A(net821),
    .B(net656),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00835_));
 sky130_fd_sc_hd__and2_1 _10205_ (.A(net825),
    .B(net660),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00836_));
 sky130_fd_sc_hd__and2_1 _10206_ (.A(net822),
    .B(net657),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00837_));
 sky130_fd_sc_hd__and2_1 _10207_ (.A(net825),
    .B(net660),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00838_));
 sky130_fd_sc_hd__and2_1 _10208_ (.A(net824),
    .B(net659),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00839_));
 sky130_fd_sc_hd__and2_1 _10209_ (.A(net824),
    .B(net659),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00840_));
 sky130_fd_sc_hd__and2_1 _10210_ (.A(net824),
    .B(net659),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00841_));
 sky130_fd_sc_hd__and2_1 _10211_ (.A(net824),
    .B(net659),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00842_));
 sky130_fd_sc_hd__and2_1 _10212_ (.A(net823),
    .B(net658),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00843_));
 sky130_fd_sc_hd__and2_1 _10213_ (.A(net823),
    .B(net658),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00844_));
 sky130_fd_sc_hd__and2_1 _10214_ (.A(net820),
    .B(net655),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00845_));
 sky130_fd_sc_hd__and2_1 _10215_ (.A(net820),
    .B(net655),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00846_));
 sky130_fd_sc_hd__and2_1 _10216_ (.A(net827),
    .B(net662),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00847_));
 sky130_fd_sc_hd__and2_1 _10217_ (.A(net827),
    .B(net662),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00848_));
 sky130_fd_sc_hd__and2_1 _10218_ (.A(net807),
    .B(net642),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00849_));
 sky130_fd_sc_hd__and2_1 _10219_ (.A(net807),
    .B(net642),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00850_));
 sky130_fd_sc_hd__and2_1 _10220_ (.A(net815),
    .B(net650),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00851_));
 sky130_fd_sc_hd__and2_1 _10221_ (.A(net815),
    .B(net650),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00852_));
 sky130_fd_sc_hd__and2_1 _10222_ (.A(net815),
    .B(net650),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00853_));
 sky130_fd_sc_hd__and2_1 _10223_ (.A(net813),
    .B(net648),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00854_));
 sky130_fd_sc_hd__and2_1 _10224_ (.A(net813),
    .B(net648),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00855_));
 sky130_fd_sc_hd__and2_1 _10225_ (.A(net813),
    .B(net648),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00856_));
 sky130_fd_sc_hd__and2_1 _10226_ (.A(net815),
    .B(net650),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00857_));
 sky130_fd_sc_hd__and2_1 _10227_ (.A(net812),
    .B(net647),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00858_));
 sky130_fd_sc_hd__and2_1 _10228_ (.A(net810),
    .B(net645),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00859_));
 sky130_fd_sc_hd__and2_1 _10229_ (.A(net810),
    .B(net645),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00860_));
 sky130_fd_sc_hd__and2_1 _10230_ (.A(net802),
    .B(net637),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00861_));
 sky130_fd_sc_hd__and2_1 _10231_ (.A(net803),
    .B(net638),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00862_));
 sky130_fd_sc_hd__and2_1 _10232_ (.A(net802),
    .B(net637),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00863_));
 sky130_fd_sc_hd__and2_1 _10233_ (.A(net803),
    .B(net638),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00864_));
 sky130_fd_sc_hd__and2_1 _10234_ (.A(net800),
    .B(net635),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00865_));
 sky130_fd_sc_hd__and2_1 _10235_ (.A(net800),
    .B(net635),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00866_));
 sky130_fd_sc_hd__and2_1 _10236_ (.A(net799),
    .B(net634),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00867_));
 sky130_fd_sc_hd__and2_1 _10237_ (.A(net804),
    .B(net639),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00868_));
 sky130_fd_sc_hd__and2_1 _10238_ (.A(net804),
    .B(net639),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00869_));
 sky130_fd_sc_hd__and2_1 _10239_ (.A(net804),
    .B(net639),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00870_));
 sky130_fd_sc_hd__and2_1 _10240_ (.A(net805),
    .B(net640),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00871_));
 sky130_fd_sc_hd__and2_1 _10241_ (.A(net805),
    .B(net640),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00872_));
 sky130_fd_sc_hd__and2_1 _10242_ (.A(net818),
    .B(net653),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00873_));
 sky130_fd_sc_hd__and2_1 _10243_ (.A(net818),
    .B(net653),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00874_));
 sky130_fd_sc_hd__and2_1 _10244_ (.A(net817),
    .B(net652),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00875_));
 sky130_fd_sc_hd__and2_1 _10245_ (.A(net818),
    .B(net653),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00876_));
 sky130_fd_sc_hd__and2_1 _10246_ (.A(net819),
    .B(net654),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00877_));
 sky130_fd_sc_hd__and2_1 _10247_ (.A(net819),
    .B(net654),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00878_));
 sky130_fd_sc_hd__and2_1 _10248_ (.A(net819),
    .B(net654),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00879_));
 sky130_fd_sc_hd__and2_1 _10249_ (.A(net753),
    .B(net588),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00880_));
 sky130_fd_sc_hd__and2_1 _10250_ (.A(net772),
    .B(net607),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00881_));
 sky130_fd_sc_hd__and2_1 _10251_ (.A(net729),
    .B(net564),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00882_));
 sky130_fd_sc_hd__and2_1 _10252_ (.A(net725),
    .B(net560),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00883_));
 sky130_fd_sc_hd__and2_1 _10253_ (.A(net725),
    .B(net560),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00884_));
 sky130_fd_sc_hd__and2_1 _10254_ (.A(net721),
    .B(net556),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00885_));
 sky130_fd_sc_hd__and2_1 _10255_ (.A(net721),
    .B(net556),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00886_));
 sky130_fd_sc_hd__and2_1 _10256_ (.A(net717),
    .B(net552),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00887_));
 sky130_fd_sc_hd__and2_1 _10257_ (.A(net717),
    .B(net552),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00888_));
 sky130_fd_sc_hd__and2_1 _10258_ (.A(net717),
    .B(net552),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00889_));
 sky130_fd_sc_hd__and2_1 _10259_ (.A(net717),
    .B(net552),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00890_));
 sky130_fd_sc_hd__and2_1 _10260_ (.A(net716),
    .B(net551),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00891_));
 sky130_fd_sc_hd__and2_1 _10261_ (.A(net716),
    .B(net551),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00892_));
 sky130_fd_sc_hd__and2_1 _10262_ (.A(net716),
    .B(net551),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00893_));
 sky130_fd_sc_hd__and2_1 _10263_ (.A(net716),
    .B(net551),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00894_));
 sky130_fd_sc_hd__and2_1 _10264_ (.A(net717),
    .B(net552),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00895_));
 sky130_fd_sc_hd__and2_1 _10265_ (.A(net717),
    .B(net552),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00896_));
 sky130_fd_sc_hd__and2_1 _10266_ (.A(net721),
    .B(net556),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00897_));
 sky130_fd_sc_hd__and2_1 _10267_ (.A(net718),
    .B(net553),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00898_));
 sky130_fd_sc_hd__and2_1 _10268_ (.A(net721),
    .B(net556),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00899_));
 sky130_fd_sc_hd__and2_1 _10269_ (.A(net723),
    .B(net558),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00900_));
 sky130_fd_sc_hd__and2_1 _10270_ (.A(net723),
    .B(net558),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00901_));
 sky130_fd_sc_hd__and2_1 _10271_ (.A(net722),
    .B(net557),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00902_));
 sky130_fd_sc_hd__and2_1 _10272_ (.A(net722),
    .B(net557),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00903_));
 sky130_fd_sc_hd__and2_1 _10273_ (.A(net722),
    .B(net557),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00904_));
 sky130_fd_sc_hd__and2_1 _10274_ (.A(net721),
    .B(net556),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00905_));
 sky130_fd_sc_hd__and2_1 _10275_ (.A(net721),
    .B(net556),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00906_));
 sky130_fd_sc_hd__and2_1 _10276_ (.A(net721),
    .B(net556),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00907_));
 sky130_fd_sc_hd__and2_1 _10277_ (.A(net721),
    .B(net556),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00908_));
 sky130_fd_sc_hd__and2_1 _10278_ (.A(net717),
    .B(net552),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00909_));
 sky130_fd_sc_hd__and2_1 _10279_ (.A(net717),
    .B(net552),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00910_));
 sky130_fd_sc_hd__and2_1 _10280_ (.A(net717),
    .B(net552),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00911_));
 sky130_fd_sc_hd__and2_1 _10281_ (.A(net716),
    .B(net551),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00912_));
 sky130_fd_sc_hd__and2_1 _10282_ (.A(net716),
    .B(net551),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00913_));
 sky130_fd_sc_hd__and2_1 _10283_ (.A(net716),
    .B(net551),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00914_));
 sky130_fd_sc_hd__and2_1 _10284_ (.A(net833),
    .B(net668),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00915_));
 sky130_fd_sc_hd__and2_1 _10285_ (.A(net828),
    .B(net663),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00916_));
 sky130_fd_sc_hd__and2_1 _10286_ (.A(net828),
    .B(net663),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00917_));
 sky130_fd_sc_hd__and2_1 _10287_ (.A(net831),
    .B(net666),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00918_));
 sky130_fd_sc_hd__and2_1 _10288_ (.A(net833),
    .B(net668),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00919_));
 sky130_fd_sc_hd__and2_1 _10289_ (.A(net833),
    .B(net668),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00920_));
 sky130_fd_sc_hd__and2_1 _10290_ (.A(net829),
    .B(net664),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00921_));
 sky130_fd_sc_hd__and2_1 _10291_ (.A(net829),
    .B(net664),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00922_));
 sky130_fd_sc_hd__and2_1 _10292_ (.A(net857),
    .B(net692),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00923_));
 sky130_fd_sc_hd__and2_1 _10293_ (.A(net861),
    .B(net696),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00924_));
 sky130_fd_sc_hd__and2_1 _10294_ (.A(net829),
    .B(net664),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00925_));
 sky130_fd_sc_hd__and2_1 _10295_ (.A(net861),
    .B(net696),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00926_));
 sky130_fd_sc_hd__and2_1 _10296_ (.A(net859),
    .B(net694),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00927_));
 sky130_fd_sc_hd__and2_1 _10297_ (.A(net859),
    .B(net694),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00928_));
 sky130_fd_sc_hd__and2_1 _10298_ (.A(net859),
    .B(net694),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00929_));
 sky130_fd_sc_hd__and2_1 _10299_ (.A(net857),
    .B(net692),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00930_));
 sky130_fd_sc_hd__and2_1 _10300_ (.A(net855),
    .B(net690),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00931_));
 sky130_fd_sc_hd__and2_1 _10301_ (.A(net856),
    .B(net691),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00932_));
 sky130_fd_sc_hd__and2_1 _10302_ (.A(net843),
    .B(net678),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00933_));
 sky130_fd_sc_hd__and2_1 _10303_ (.A(net844),
    .B(net679),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00934_));
 sky130_fd_sc_hd__and2_1 _10304_ (.A(net844),
    .B(net679),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00935_));
 sky130_fd_sc_hd__and2_1 _10305_ (.A(net841),
    .B(net676),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00936_));
 sky130_fd_sc_hd__and2_1 _10306_ (.A(net840),
    .B(net675),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00937_));
 sky130_fd_sc_hd__and2_1 _10307_ (.A(net840),
    .B(net675),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00938_));
 sky130_fd_sc_hd__and2_1 _10308_ (.A(net839),
    .B(net674),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00939_));
 sky130_fd_sc_hd__and2_1 _10309_ (.A(net839),
    .B(net674),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00940_));
 sky130_fd_sc_hd__and2_1 _10310_ (.A(net839),
    .B(net674),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00941_));
 sky130_fd_sc_hd__and2_1 _10311_ (.A(net838),
    .B(net673),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00942_));
 sky130_fd_sc_hd__and2_1 _10312_ (.A(net785),
    .B(net620),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00943_));
 sky130_fd_sc_hd__and2_1 _10313_ (.A(net784),
    .B(net619),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00944_));
 sky130_fd_sc_hd__and2_1 _10314_ (.A(net784),
    .B(net619),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00945_));
 sky130_fd_sc_hd__and2_1 _10315_ (.A(net779),
    .B(net614),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00946_));
 sky130_fd_sc_hd__and2_1 _10316_ (.A(net731),
    .B(net566),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00947_));
 sky130_fd_sc_hd__and2_1 _10317_ (.A(net758),
    .B(net593),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00948_));
 sky130_fd_sc_hd__and2_1 _10318_ (.A(net758),
    .B(net593),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00949_));
 sky130_fd_sc_hd__and2_1 _10319_ (.A(net758),
    .B(net593),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00950_));
 sky130_fd_sc_hd__and2_1 _10320_ (.A(net758),
    .B(net593),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00951_));
 sky130_fd_sc_hd__and2_1 _10321_ (.A(net758),
    .B(net593),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00952_));
 sky130_fd_sc_hd__and2_1 _10322_ (.A(net730),
    .B(net565),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00953_));
 sky130_fd_sc_hd__and2_1 _10323_ (.A(net730),
    .B(net565),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00954_));
 sky130_fd_sc_hd__and2_1 _10324_ (.A(net731),
    .B(net566),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00955_));
 sky130_fd_sc_hd__and2_1 _10325_ (.A(net728),
    .B(net563),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00956_));
 sky130_fd_sc_hd__and2_1 _10326_ (.A(net728),
    .B(net563),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00957_));
 sky130_fd_sc_hd__and2_1 _10327_ (.A(net730),
    .B(net565),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00958_));
 sky130_fd_sc_hd__and2_1 _10328_ (.A(net767),
    .B(net602),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00959_));
 sky130_fd_sc_hd__and2_1 _10329_ (.A(net768),
    .B(net603),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00960_));
 sky130_fd_sc_hd__and2_1 _10330_ (.A(net767),
    .B(net602),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00961_));
 sky130_fd_sc_hd__and2_1 _10331_ (.A(net728),
    .B(net563),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00962_));
 sky130_fd_sc_hd__and2_1 _10332_ (.A(net774),
    .B(net609),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00963_));
 sky130_fd_sc_hd__and2_1 _10333_ (.A(net767),
    .B(net602),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00964_));
 sky130_fd_sc_hd__and2_1 _10334_ (.A(net774),
    .B(net609),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00965_));
 sky130_fd_sc_hd__and2_1 _10335_ (.A(net768),
    .B(net603),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00966_));
 sky130_fd_sc_hd__and2_1 _10336_ (.A(net768),
    .B(net603),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00967_));
 sky130_fd_sc_hd__and2_1 _10337_ (.A(net728),
    .B(net563),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00968_));
 sky130_fd_sc_hd__and2_1 _10338_ (.A(net730),
    .B(net565),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00969_));
 sky130_fd_sc_hd__and2_1 _10339_ (.A(net727),
    .B(net562),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00970_));
 sky130_fd_sc_hd__and2_1 _10340_ (.A(net768),
    .B(net603),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00971_));
 sky130_fd_sc_hd__and2_1 _10341_ (.A(net727),
    .B(net562),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00972_));
 sky130_fd_sc_hd__and2_1 _10342_ (.A(net729),
    .B(net564),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00973_));
 sky130_fd_sc_hd__and2_1 _10343_ (.A(net775),
    .B(net610),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00974_));
 sky130_fd_sc_hd__and2_1 _10344_ (.A(net775),
    .B(net610),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00975_));
 sky130_fd_sc_hd__and2_1 _10345_ (.A(net776),
    .B(net611),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00976_));
 sky130_fd_sc_hd__and2_1 _10346_ (.A(net776),
    .B(net611),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00977_));
 sky130_fd_sc_hd__and2_1 _10347_ (.A(net774),
    .B(net609),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00978_));
 sky130_fd_sc_hd__and2_1 _10348_ (.A(net775),
    .B(net610),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00979_));
 sky130_fd_sc_hd__and2_1 _10349_ (.A(net775),
    .B(net610),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00980_));
 sky130_fd_sc_hd__and2_1 _10350_ (.A(net774),
    .B(net609),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00981_));
 sky130_fd_sc_hd__and2_1 _10351_ (.A(net729),
    .B(net564),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00982_));
 sky130_fd_sc_hd__and2_1 _10352_ (.A(net719),
    .B(net554),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00983_));
 sky130_fd_sc_hd__and2_1 _10353_ (.A(net727),
    .B(net562),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00984_));
 sky130_fd_sc_hd__and2_1 _10354_ (.A(net719),
    .B(net554),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00985_));
 sky130_fd_sc_hd__and2_1 _10355_ (.A(net727),
    .B(net562),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00986_));
 sky130_fd_sc_hd__and2_1 _10356_ (.A(net716),
    .B(net551),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00987_));
 sky130_fd_sc_hd__and2_1 _10357_ (.A(net718),
    .B(net553),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00988_));
 sky130_fd_sc_hd__and2_1 _10358_ (.A(net720),
    .B(net555),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00989_));
 sky130_fd_sc_hd__and2_1 _10359_ (.A(net716),
    .B(net551),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00990_));
 sky130_fd_sc_hd__and2_1 _10360_ (.A(net727),
    .B(net562),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00991_));
 sky130_fd_sc_hd__and2_1 _10361_ (.A(net716),
    .B(net551),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00992_));
 sky130_fd_sc_hd__and2_1 _10362_ (.A(net727),
    .B(net562),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00993_));
 sky130_fd_sc_hd__and2_1 _10363_ (.A(net718),
    .B(net553),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00994_));
 sky130_fd_sc_hd__and2_1 _10364_ (.A(net718),
    .B(net553),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00995_));
 sky130_fd_sc_hd__and2_1 _10365_ (.A(net720),
    .B(net555),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00996_));
 sky130_fd_sc_hd__and2_1 _10366_ (.A(net732),
    .B(net567),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00997_));
 sky130_fd_sc_hd__and2_1 _10367_ (.A(net758),
    .B(net593),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00998_));
 sky130_fd_sc_hd__and2_1 _10368_ (.A(net758),
    .B(net593),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00999_));
 sky130_fd_sc_hd__and2_1 _10369_ (.A(net758),
    .B(net593),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01000_));
 sky130_fd_sc_hd__and2_1 _10370_ (.A(net758),
    .B(net593),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01001_));
 sky130_fd_sc_hd__and2_1 _10371_ (.A(net760),
    .B(net595),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01002_));
 sky130_fd_sc_hd__and2_1 _10372_ (.A(net760),
    .B(net595),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01003_));
 sky130_fd_sc_hd__and2_1 _10373_ (.A(net760),
    .B(net595),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01004_));
 sky130_fd_sc_hd__and2_1 _10374_ (.A(net760),
    .B(net595),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01005_));
 sky130_fd_sc_hd__and2_1 _10375_ (.A(net761),
    .B(net596),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01006_));
 sky130_fd_sc_hd__and2_1 _10376_ (.A(net761),
    .B(net596),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01007_));
 sky130_fd_sc_hd__and2_1 _10377_ (.A(net759),
    .B(net594),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01008_));
 sky130_fd_sc_hd__and2_1 _10378_ (.A(net759),
    .B(net594),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01009_));
 sky130_fd_sc_hd__and2_1 _10379_ (.A(net769),
    .B(net604),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01010_));
 sky130_fd_sc_hd__and2_1 _10380_ (.A(net769),
    .B(net604),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01011_));
 sky130_fd_sc_hd__and2_1 _10381_ (.A(net769),
    .B(net604),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01012_));
 sky130_fd_sc_hd__and2_1 _10382_ (.A(net769),
    .B(net604),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01013_));
 sky130_fd_sc_hd__and2_1 _10383_ (.A(net762),
    .B(net597),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01014_));
 sky130_fd_sc_hd__and2_1 _10384_ (.A(net760),
    .B(net595),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01015_));
 sky130_fd_sc_hd__and2_1 _10385_ (.A(net762),
    .B(net597),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01016_));
 sky130_fd_sc_hd__and2_1 _10386_ (.A(net762),
    .B(net597),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01017_));
 sky130_fd_sc_hd__and2_1 _10387_ (.A(net769),
    .B(net604),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01018_));
 sky130_fd_sc_hd__and2_1 _10388_ (.A(net769),
    .B(net604),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01019_));
 sky130_fd_sc_hd__and2_1 _10389_ (.A(net770),
    .B(net605),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01020_));
 sky130_fd_sc_hd__and2_1 _10390_ (.A(net769),
    .B(net604),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01021_));
 sky130_fd_sc_hd__and2_1 _10391_ (.A(net735),
    .B(net570),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01022_));
 sky130_fd_sc_hd__and2_1 _10392_ (.A(net748),
    .B(net583),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01023_));
 sky130_fd_sc_hd__and2_1 _10393_ (.A(net748),
    .B(net583),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01024_));
 sky130_fd_sc_hd__and2_1 _10394_ (.A(net801),
    .B(net636),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01025_));
 sky130_fd_sc_hd__and2_1 _10395_ (.A(net801),
    .B(net636),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01026_));
 sky130_fd_sc_hd__and2_1 _10396_ (.A(net801),
    .B(net636),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01027_));
 sky130_fd_sc_hd__and2_1 _10397_ (.A(net801),
    .B(net636),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01028_));
 sky130_fd_sc_hd__and2_1 _10398_ (.A(net801),
    .B(net636),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01029_));
 sky130_fd_sc_hd__and2_1 _10399_ (.A(net801),
    .B(net636),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01030_));
 sky130_fd_sc_hd__and2_1 _10400_ (.A(net746),
    .B(net581),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01031_));
 sky130_fd_sc_hd__and2_1 _10401_ (.A(net746),
    .B(net581),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01032_));
 sky130_fd_sc_hd__and2_1 _10402_ (.A(net747),
    .B(net582),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01033_));
 sky130_fd_sc_hd__and2_1 _10403_ (.A(net747),
    .B(net582),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01034_));
 sky130_fd_sc_hd__and2_1 _10404_ (.A(net746),
    .B(net581),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01035_));
 sky130_fd_sc_hd__and2_1 _10405_ (.A(net746),
    .B(net581),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01036_));
 sky130_fd_sc_hd__and2_1 _10406_ (.A(net746),
    .B(net581),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01037_));
 sky130_fd_sc_hd__and2_1 _10407_ (.A(net746),
    .B(net581),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01038_));
 sky130_fd_sc_hd__and2_1 _10408_ (.A(net741),
    .B(net576),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01039_));
 sky130_fd_sc_hd__and2_1 _10409_ (.A(net742),
    .B(net577),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01040_));
 sky130_fd_sc_hd__and2_1 _10410_ (.A(net738),
    .B(net573),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01041_));
 sky130_fd_sc_hd__and2_1 _10411_ (.A(net741),
    .B(net576),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01042_));
 sky130_fd_sc_hd__and2_1 _10412_ (.A(net739),
    .B(net574),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01043_));
 sky130_fd_sc_hd__and2_1 _10413_ (.A(net742),
    .B(net577),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01044_));
 sky130_fd_sc_hd__and2_1 _10414_ (.A(net737),
    .B(net572),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01045_));
 sky130_fd_sc_hd__and2_1 _10415_ (.A(net742),
    .B(net577),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01046_));
 sky130_fd_sc_hd__and2_1 _10416_ (.A(net737),
    .B(net572),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01047_));
 sky130_fd_sc_hd__and2_1 _10417_ (.A(net740),
    .B(net575),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01048_));
 sky130_fd_sc_hd__and2_1 _10418_ (.A(net740),
    .B(net575),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01049_));
 sky130_fd_sc_hd__and2_1 _10419_ (.A(net740),
    .B(net575),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01050_));
 sky130_fd_sc_hd__and2_1 _10420_ (.A(net739),
    .B(net574),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01051_));
 sky130_fd_sc_hd__and2_1 _10421_ (.A(net739),
    .B(net574),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01052_));
 sky130_fd_sc_hd__and2_1 _10422_ (.A(net739),
    .B(net574),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01053_));
 sky130_fd_sc_hd__and2_1 _10423_ (.A(net739),
    .B(net574),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01054_));
 sky130_fd_sc_hd__and2_1 _10424_ (.A(net763),
    .B(net598),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01055_));
 sky130_fd_sc_hd__and2_1 _10425_ (.A(net766),
    .B(net601),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01056_));
 sky130_fd_sc_hd__and2_1 _10426_ (.A(net821),
    .B(net656),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01057_));
 sky130_fd_sc_hd__and2_1 _10427_ (.A(net818),
    .B(net653),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01058_));
 sky130_fd_sc_hd__and2_1 _10428_ (.A(net818),
    .B(net653),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01059_));
 sky130_fd_sc_hd__and2_1 _10429_ (.A(net818),
    .B(net653),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01060_));
 sky130_fd_sc_hd__and2_1 _10430_ (.A(net822),
    .B(net657),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01061_));
 sky130_fd_sc_hd__and2_1 _10431_ (.A(net822),
    .B(net657),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01062_));
 sky130_fd_sc_hd__and2_1 _10432_ (.A(net822),
    .B(net657),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01063_));
 sky130_fd_sc_hd__and2_1 _10433_ (.A(net823),
    .B(net658),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01064_));
 sky130_fd_sc_hd__and2_1 _10434_ (.A(net820),
    .B(net655),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01065_));
 sky130_fd_sc_hd__and2_1 _10435_ (.A(net820),
    .B(net655),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01066_));
 sky130_fd_sc_hd__and2_1 _10436_ (.A(net818),
    .B(net653),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01067_));
 sky130_fd_sc_hd__and2_1 _10437_ (.A(net820),
    .B(net655),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01068_));
 sky130_fd_sc_hd__and2_1 _10438_ (.A(net820),
    .B(net655),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01069_));
 sky130_fd_sc_hd__and2_1 _10439_ (.A(net819),
    .B(net654),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01070_));
 sky130_fd_sc_hd__and2_1 _10440_ (.A(net827),
    .B(net662),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01071_));
 sky130_fd_sc_hd__and2_1 _10441_ (.A(net819),
    .B(net654),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01072_));
 sky130_fd_sc_hd__and2_1 _10442_ (.A(net807),
    .B(net642),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01073_));
 sky130_fd_sc_hd__and2_1 _10443_ (.A(net807),
    .B(net642),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01074_));
 sky130_fd_sc_hd__and2_1 _10444_ (.A(net806),
    .B(net641),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01075_));
 sky130_fd_sc_hd__and2_1 _10445_ (.A(net806),
    .B(net641),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01076_));
 sky130_fd_sc_hd__and2_1 _10446_ (.A(net815),
    .B(net650),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01077_));
 sky130_fd_sc_hd__and2_1 _10447_ (.A(net815),
    .B(net650),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01078_));
 sky130_fd_sc_hd__and2_1 _10448_ (.A(net813),
    .B(net648),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01079_));
 sky130_fd_sc_hd__and2_1 _10449_ (.A(net813),
    .B(net648),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01080_));
 sky130_fd_sc_hd__and2_1 _10450_ (.A(net810),
    .B(net645),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01081_));
 sky130_fd_sc_hd__and2_1 _10451_ (.A(net812),
    .B(net647),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01082_));
 sky130_fd_sc_hd__and2_1 _10452_ (.A(net809),
    .B(net644),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01083_));
 sky130_fd_sc_hd__and2_1 _10453_ (.A(net809),
    .B(net644),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01084_));
 sky130_fd_sc_hd__and2_1 _10454_ (.A(net803),
    .B(net638),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01085_));
 sky130_fd_sc_hd__and2_1 _10455_ (.A(net802),
    .B(net637),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01086_));
 sky130_fd_sc_hd__and2_1 _10456_ (.A(net802),
    .B(net637),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01087_));
 sky130_fd_sc_hd__and2_1 _10457_ (.A(net803),
    .B(net638),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01088_));
 sky130_fd_sc_hd__and2_1 _10458_ (.A(net735),
    .B(net570),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01089_));
 sky130_fd_sc_hd__and2_1 _10459_ (.A(net735),
    .B(net570),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01090_));
 sky130_fd_sc_hd__and2_1 _10460_ (.A(net766),
    .B(net601),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01091_));
 sky130_fd_sc_hd__and2_1 _10461_ (.A(net828),
    .B(net663),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01092_));
 sky130_fd_sc_hd__and2_1 _10462_ (.A(net828),
    .B(net663),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01093_));
 sky130_fd_sc_hd__and2_1 _10463_ (.A(net828),
    .B(net663),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01094_));
 sky130_fd_sc_hd__and2_1 _10464_ (.A(net828),
    .B(net663),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01095_));
 sky130_fd_sc_hd__and2_1 _10465_ (.A(net828),
    .B(net663),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01096_));
 sky130_fd_sc_hd__and2_1 _10466_ (.A(net829),
    .B(net664),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01097_));
 sky130_fd_sc_hd__and2_1 _10467_ (.A(net829),
    .B(net664),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01098_));
 sky130_fd_sc_hd__and2_1 _10468_ (.A(net829),
    .B(net664),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01099_));
 sky130_fd_sc_hd__and2_1 _10469_ (.A(net829),
    .B(net664),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01100_));
 sky130_fd_sc_hd__and2_1 _10470_ (.A(net829),
    .B(net664),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01101_));
 sky130_fd_sc_hd__and2_1 _10471_ (.A(net830),
    .B(net665),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01102_));
 sky130_fd_sc_hd__and2_1 _10472_ (.A(net830),
    .B(net665),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01103_));
 sky130_fd_sc_hd__and2_1 _10473_ (.A(net855),
    .B(net690),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01104_));
 sky130_fd_sc_hd__and2_1 _10474_ (.A(net855),
    .B(net690),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01105_));
 sky130_fd_sc_hd__and2_1 _10475_ (.A(net855),
    .B(net690),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01106_));
 sky130_fd_sc_hd__and2_1 _10476_ (.A(net856),
    .B(net691),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01107_));
 sky130_fd_sc_hd__and2_1 _10477_ (.A(net841),
    .B(net676),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01108_));
 sky130_fd_sc_hd__and2_1 _10478_ (.A(net841),
    .B(net676),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01109_));
 sky130_fd_sc_hd__and2_1 _10479_ (.A(net841),
    .B(net676),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01110_));
 sky130_fd_sc_hd__and2_1 _10480_ (.A(net840),
    .B(net675),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01111_));
 sky130_fd_sc_hd__and2_1 _10481_ (.A(net840),
    .B(net675),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01112_));
 sky130_fd_sc_hd__and2_1 _10482_ (.A(net840),
    .B(net675),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01113_));
 sky130_fd_sc_hd__and2_1 _10483_ (.A(net840),
    .B(net675),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01114_));
 sky130_fd_sc_hd__and2_1 _10484_ (.A(net837),
    .B(net672),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01115_));
 sky130_fd_sc_hd__and2_1 _10485_ (.A(net839),
    .B(net674),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01116_));
 sky130_fd_sc_hd__and2_1 _10486_ (.A(net839),
    .B(net674),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01117_));
 sky130_fd_sc_hd__and2_1 _10487_ (.A(net838),
    .B(net673),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01118_));
 sky130_fd_sc_hd__and2_1 _10488_ (.A(net785),
    .B(net620),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01119_));
 sky130_fd_sc_hd__and2_1 _10489_ (.A(net785),
    .B(net620),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01120_));
 sky130_fd_sc_hd__and2_1 _10490_ (.A(net779),
    .B(net614),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01121_));
 sky130_fd_sc_hd__and2_1 _10491_ (.A(net779),
    .B(net614),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01122_));
 sky130_fd_sc_hd__and2_1 _10492_ (.A(net780),
    .B(net615),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01123_));
 sky130_fd_sc_hd__and2_1 _10493_ (.A(net753),
    .B(net588),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01124_));
 sky130_fd_sc_hd__and2_1 _10494_ (.A(net752),
    .B(net587),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01125_));
 sky130_fd_sc_hd__and2_1 _10495_ (.A(net732),
    .B(net567),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01126_));
 sky130_fd_sc_hd__and2_1 _10496_ (.A(net755),
    .B(net590),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01127_));
 sky130_fd_sc_hd__and2_1 _10497_ (.A(net755),
    .B(net590),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01128_));
 sky130_fd_sc_hd__and2_1 _10498_ (.A(net751),
    .B(net586),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01129_));
 sky130_fd_sc_hd__and2_1 _10499_ (.A(net755),
    .B(net590),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01130_));
 sky130_fd_sc_hd__and2_1 _10500_ (.A(net734),
    .B(net569),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01131_));
 sky130_fd_sc_hd__and2_1 _10501_ (.A(net734),
    .B(net569),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01132_));
 sky130_fd_sc_hd__and2_1 _10502_ (.A(net734),
    .B(net569),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01133_));
 sky130_fd_sc_hd__and2_1 _10503_ (.A(net730),
    .B(net565),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01134_));
 sky130_fd_sc_hd__and2_1 _10504_ (.A(net750),
    .B(net585),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01135_));
 sky130_fd_sc_hd__and2_1 _10505_ (.A(net750),
    .B(net585),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01136_));
 sky130_fd_sc_hd__and2_1 _10506_ (.A(net750),
    .B(net585),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01137_));
 sky130_fd_sc_hd__and2_1 _10507_ (.A(net754),
    .B(net589),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01138_));
 sky130_fd_sc_hd__and2_1 _10508_ (.A(net754),
    .B(net589),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01139_));
 sky130_fd_sc_hd__and2_1 _10509_ (.A(net754),
    .B(net589),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01140_));
 sky130_fd_sc_hd__and2_1 _10510_ (.A(net757),
    .B(net592),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01141_));
 sky130_fd_sc_hd__and2_1 _10511_ (.A(net757),
    .B(net592),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01142_));
 sky130_fd_sc_hd__and2_1 _10512_ (.A(net757),
    .B(net592),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01143_));
 sky130_fd_sc_hd__and2_1 _10513_ (.A(net755),
    .B(net590),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01144_));
 sky130_fd_sc_hd__and2_1 _10514_ (.A(net756),
    .B(net591),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01145_));
 sky130_fd_sc_hd__and2_1 _10515_ (.A(net756),
    .B(net591),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01146_));
 sky130_fd_sc_hd__and2_1 _10516_ (.A(net755),
    .B(net590),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01147_));
 sky130_fd_sc_hd__and2_1 _10517_ (.A(net755),
    .B(net590),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01148_));
 sky130_fd_sc_hd__and2_1 _10518_ (.A(net733),
    .B(net568),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01149_));
 sky130_fd_sc_hd__and2_1 _10519_ (.A(net733),
    .B(net568),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01150_));
 sky130_fd_sc_hd__and2_1 _10520_ (.A(net734),
    .B(net569),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01151_));
 sky130_fd_sc_hd__and2_1 _10521_ (.A(net733),
    .B(net568),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01152_));
 sky130_fd_sc_hd__and2_1 _10522_ (.A(net733),
    .B(net568),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01153_));
 sky130_fd_sc_hd__and2_1 _10523_ (.A(net725),
    .B(net560),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01154_));
 sky130_fd_sc_hd__and2_1 _10524_ (.A(net800),
    .B(net635),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01155_));
 sky130_fd_sc_hd__and2_1 _10525_ (.A(net799),
    .B(net634),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01156_));
 sky130_fd_sc_hd__and2_1 _10526_ (.A(net799),
    .B(net634),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01157_));
 sky130_fd_sc_hd__and2_1 _10527_ (.A(net804),
    .B(net639),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01158_));
 sky130_fd_sc_hd__and2_1 _10528_ (.A(net804),
    .B(net639),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01159_));
 sky130_fd_sc_hd__and2_1 _10529_ (.A(net805),
    .B(net640),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01160_));
 sky130_fd_sc_hd__and2_1 _10530_ (.A(net805),
    .B(net640),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01161_));
 sky130_fd_sc_hd__and2_1 _10531_ (.A(net805),
    .B(net640),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01162_));
 sky130_fd_sc_hd__and2_1 _10532_ (.A(net817),
    .B(net652),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01163_));
 sky130_fd_sc_hd__and2_1 _10533_ (.A(net817),
    .B(net652),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01164_));
 sky130_fd_sc_hd__and2_1 _10534_ (.A(net817),
    .B(net652),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01165_));
 sky130_fd_sc_hd__and2_1 _10535_ (.A(net817),
    .B(net652),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01166_));
 sky130_fd_sc_hd__and2_1 _10536_ (.A(net817),
    .B(net652),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01167_));
 sky130_fd_sc_hd__and2_1 _10537_ (.A(net819),
    .B(net654),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01168_));
 sky130_fd_sc_hd__and2_1 _10538_ (.A(net717),
    .B(net552),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01169_));
 sky130_fd_sc_hd__and2_1 _10539_ (.A(net728),
    .B(net563),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01170_));
 sky130_fd_sc_hd__and2_1 _10540_ (.A(net731),
    .B(net566),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01171_));
 sky130_fd_sc_hd__and2_1 _10541_ (.A(net730),
    .B(net565),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01172_));
 sky130_fd_sc_hd__and2_1 _10542_ (.A(net731),
    .B(net566),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01173_));
 sky130_fd_sc_hd__and2_1 _10543_ (.A(net730),
    .B(net565),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01174_));
 sky130_fd_sc_hd__and2_1 _10544_ (.A(net728),
    .B(net563),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01175_));
 sky130_fd_sc_hd__and2_1 _10545_ (.A(net736),
    .B(net571),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01176_));
 sky130_fd_sc_hd__and2_1 _10546_ (.A(net833),
    .B(net668),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01177_));
 sky130_fd_sc_hd__and2_1 _10547_ (.A(net832),
    .B(net667),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01178_));
 sky130_fd_sc_hd__and2_1 _10548_ (.A(net834),
    .B(net669),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01179_));
 sky130_fd_sc_hd__and2_1 _10549_ (.A(net834),
    .B(net669),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01180_));
 sky130_fd_sc_hd__and2_1 _10550_ (.A(net832),
    .B(net667),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01181_));
 sky130_fd_sc_hd__and2_1 _10551_ (.A(net832),
    .B(net667),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01182_));
 sky130_fd_sc_hd__and2_1 _10552_ (.A(net832),
    .B(net667),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01183_));
 sky130_fd_sc_hd__and2_1 _10553_ (.A(net832),
    .B(net667),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01184_));
 sky130_fd_sc_hd__and2_1 _10554_ (.A(net862),
    .B(net697),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01185_));
 sky130_fd_sc_hd__and2_1 _10555_ (.A(net834),
    .B(net669),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01186_));
 sky130_fd_sc_hd__and2_1 _10556_ (.A(net834),
    .B(net669),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01187_));
 sky130_fd_sc_hd__and2_1 _10557_ (.A(net860),
    .B(net695),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01188_));
 sky130_fd_sc_hd__and2_1 _10558_ (.A(net860),
    .B(net695),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01189_));
 sky130_fd_sc_hd__and2_1 _10559_ (.A(net860),
    .B(net695),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01190_));
 sky130_fd_sc_hd__and2_1 _10560_ (.A(net862),
    .B(net697),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01191_));
 sky130_fd_sc_hd__and2_1 _10561_ (.A(net862),
    .B(net697),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01192_));
 sky130_fd_sc_hd__and2_1 _10562_ (.A(net860),
    .B(net695),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01193_));
 sky130_fd_sc_hd__and2_1 _10563_ (.A(net861),
    .B(net696),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01194_));
 sky130_fd_sc_hd__and2_1 _10564_ (.A(net862),
    .B(net697),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01195_));
 sky130_fd_sc_hd__and2_1 _10565_ (.A(net862),
    .B(net697),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01196_));
 sky130_fd_sc_hd__and2_1 _10566_ (.A(net864),
    .B(net699),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01197_));
 sky130_fd_sc_hd__and2_1 _10567_ (.A(net862),
    .B(net697),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01198_));
 sky130_fd_sc_hd__and2_1 _10568_ (.A(net861),
    .B(net696),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01199_));
 sky130_fd_sc_hd__and2_1 _10569_ (.A(net860),
    .B(net695),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01200_));
 sky130_fd_sc_hd__and2_1 _10570_ (.A(net839),
    .B(net674),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01201_));
 sky130_fd_sc_hd__and2_1 _10571_ (.A(net860),
    .B(net695),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01202_));
 sky130_fd_sc_hd__and2_1 _10572_ (.A(net860),
    .B(net695),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01203_));
 sky130_fd_sc_hd__and2_1 _10573_ (.A(net833),
    .B(net668),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01204_));
 sky130_fd_sc_hd__and2_1 _10574_ (.A(net838),
    .B(net673),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01205_));
 sky130_fd_sc_hd__and2_1 _10575_ (.A(net785),
    .B(net620),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01206_));
 sky130_fd_sc_hd__and2_1 _10576_ (.A(net784),
    .B(net619),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01207_));
 sky130_fd_sc_hd__and2_1 _10577_ (.A(net785),
    .B(net620),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01208_));
 sky130_fd_sc_hd__and2_1 _10578_ (.A(net727),
    .B(net562),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01209_));
 sky130_fd_sc_hd__and2_1 _10579_ (.A(net862),
    .B(net697),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01210_));
 sky130_fd_sc_hd__and2_1 _10580_ (.A(net799),
    .B(net634),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01211_));
 sky130_fd_sc_hd__and2_1 _10581_ (.A(net738),
    .B(net573),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01212_));
 sky130_fd_sc_hd__and2_1 _10582_ (.A(net745),
    .B(net580),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01213_));
 sky130_fd_sc_hd__and2_1 _10583_ (.A(net745),
    .B(net580),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01214_));
 sky130_fd_sc_hd__and2_1 _10584_ (.A(net797),
    .B(net632),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01215_));
 sky130_fd_sc_hd__and2_1 _10585_ (.A(net738),
    .B(net573),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01216_));
 sky130_fd_sc_hd__and2_1 _10586_ (.A(net797),
    .B(net632),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01217_));
 sky130_fd_sc_hd__and2_1 _10587_ (.A(net797),
    .B(net632),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01218_));
 sky130_fd_sc_hd__and2_1 _10588_ (.A(net738),
    .B(net573),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01219_));
 sky130_fd_sc_hd__and2_1 _10589_ (.A(net745),
    .B(net580),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01220_));
 sky130_fd_sc_hd__and2_1 _10590_ (.A(net737),
    .B(net572),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01221_));
 sky130_fd_sc_hd__and2_1 _10591_ (.A(net799),
    .B(net634),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01222_));
 sky130_fd_sc_hd__and2_1 _10592_ (.A(net799),
    .B(net634),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01223_));
 sky130_fd_sc_hd__and2_1 _10593_ (.A(net745),
    .B(net580),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01224_));
 sky130_fd_sc_hd__and2_1 _10594_ (.A(net737),
    .B(net572),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01225_));
 sky130_fd_sc_hd__and2_1 _10595_ (.A(net797),
    .B(net632),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01226_));
 sky130_fd_sc_hd__and2_1 _10596_ (.A(net797),
    .B(net632),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01227_));
 sky130_fd_sc_hd__and2_1 _10597_ (.A(net745),
    .B(net580),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01228_));
 sky130_fd_sc_hd__and2_1 _10598_ (.A(net743),
    .B(net578),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01229_));
 sky130_fd_sc_hd__and2_1 _10599_ (.A(net738),
    .B(net573),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01230_));
 sky130_fd_sc_hd__and2_1 _10600_ (.A(net799),
    .B(net634),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01231_));
 sky130_fd_sc_hd__and2_1 _10601_ (.A(net738),
    .B(net573),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01232_));
 sky130_fd_sc_hd__and2_1 _10602_ (.A(net743),
    .B(net578),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01233_));
 sky130_fd_sc_hd__and2_1 _10603_ (.A(net743),
    .B(net578),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01234_));
 sky130_fd_sc_hd__and2_1 _10604_ (.A(net738),
    .B(net573),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01235_));
 sky130_fd_sc_hd__and2_1 _10605_ (.A(net743),
    .B(net578),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01236_));
 sky130_fd_sc_hd__and2_1 _10606_ (.A(net743),
    .B(net578),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01237_));
 sky130_fd_sc_hd__and2_1 _10607_ (.A(net743),
    .B(net578),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01238_));
 sky130_fd_sc_hd__and2_1 _10608_ (.A(net745),
    .B(net580),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01239_));
 sky130_fd_sc_hd__and2_1 _10609_ (.A(net797),
    .B(net632),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01240_));
 sky130_fd_sc_hd__and2_1 _10610_ (.A(net738),
    .B(net573),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01241_));
 sky130_fd_sc_hd__and2_1 _10611_ (.A(net743),
    .B(net578),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01242_));
 sky130_fd_sc_hd__and2_1 _10612_ (.A(net771),
    .B(net606),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01243_));
 sky130_fd_sc_hd__and2_1 _10613_ (.A(net719),
    .B(net554),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01244_));
 sky130_fd_sc_hd__and2_1 _10614_ (.A(net719),
    .B(net554),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01245_));
 sky130_fd_sc_hd__and2_1 _10615_ (.A(net719),
    .B(net554),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01246_));
 sky130_fd_sc_hd__and2_1 _10616_ (.A(net718),
    .B(net553),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01247_));
 sky130_fd_sc_hd__dfxtp_1 _10617_ (.CLK(clknet_leaf_83_clk),
    .D(_01248_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _10618_ (.CLK(clknet_leaf_83_clk),
    .D(_01249_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _10619_ (.CLK(clknet_leaf_83_clk),
    .D(_01250_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _10620_ (.CLK(clknet_leaf_83_clk),
    .D(_01251_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _10621_ (.CLK(clknet_leaf_83_clk),
    .D(_01252_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _10622_ (.CLK(clknet_leaf_83_clk),
    .D(_01253_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _10623_ (.CLK(clknet_leaf_81_clk),
    .D(_01254_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 _10624_ (.CLK(clknet_leaf_82_clk),
    .D(_01255_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 _10625_ (.CLK(clknet_leaf_65_clk),
    .D(_01256_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[8] ));
 sky130_fd_sc_hd__dfxtp_1 _10626_ (.CLK(clknet_leaf_67_clk),
    .D(_01257_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[9] ));
 sky130_fd_sc_hd__dfxtp_1 _10627_ (.CLK(clknet_leaf_82_clk),
    .D(_01258_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[10] ));
 sky130_fd_sc_hd__dfxtp_1 _10628_ (.CLK(clknet_leaf_67_clk),
    .D(_01259_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[11] ));
 sky130_fd_sc_hd__dfxtp_1 _10629_ (.CLK(clknet_leaf_66_clk),
    .D(_01260_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[12] ));
 sky130_fd_sc_hd__dfxtp_1 _10630_ (.CLK(clknet_leaf_67_clk),
    .D(_01261_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[13] ));
 sky130_fd_sc_hd__dfxtp_1 _10631_ (.CLK(clknet_leaf_66_clk),
    .D(_01262_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[14] ));
 sky130_fd_sc_hd__dfxtp_1 _10632_ (.CLK(clknet_leaf_64_clk),
    .D(_01263_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[15] ));
 sky130_fd_sc_hd__dfxtp_1 _10633_ (.CLK(clknet_leaf_69_clk),
    .D(_01264_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[16] ));
 sky130_fd_sc_hd__dfxtp_1 _10634_ (.CLK(clknet_leaf_73_clk),
    .D(_01265_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[17] ));
 sky130_fd_sc_hd__dfxtp_1 _10635_ (.CLK(clknet_leaf_69_clk),
    .D(_01266_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[18] ));
 sky130_fd_sc_hd__dfxtp_1 _10636_ (.CLK(clknet_leaf_73_clk),
    .D(_01267_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[19] ));
 sky130_fd_sc_hd__dfxtp_1 _10637_ (.CLK(clknet_leaf_77_clk),
    .D(_01268_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[20] ));
 sky130_fd_sc_hd__dfxtp_1 _10638_ (.CLK(clknet_leaf_72_clk),
    .D(_01269_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[21] ));
 sky130_fd_sc_hd__dfxtp_1 _10639_ (.CLK(clknet_leaf_74_clk),
    .D(_01270_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[22] ));
 sky130_fd_sc_hd__dfxtp_1 _10640_ (.CLK(clknet_leaf_73_clk),
    .D(_01271_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[23] ));
 sky130_fd_sc_hd__dfxtp_1 _10641_ (.CLK(clknet_leaf_76_clk),
    .D(_01272_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[24] ));
 sky130_fd_sc_hd__dfxtp_1 _10642_ (.CLK(clknet_leaf_74_clk),
    .D(_01273_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[25] ));
 sky130_fd_sc_hd__dfxtp_1 _10643_ (.CLK(clknet_leaf_74_clk),
    .D(_01274_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[26] ));
 sky130_fd_sc_hd__dfxtp_1 _10644_ (.CLK(clknet_leaf_75_clk),
    .D(_01275_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[27] ));
 sky130_fd_sc_hd__dfxtp_1 _10645_ (.CLK(clknet_leaf_104_clk),
    .D(_01276_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[28] ));
 sky130_fd_sc_hd__dfxtp_1 _10646_ (.CLK(clknet_leaf_103_clk),
    .D(_01277_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[29] ));
 sky130_fd_sc_hd__dfxtp_1 _10647_ (.CLK(clknet_leaf_103_clk),
    .D(_01278_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[30] ));
 sky130_fd_sc_hd__dfxtp_1 _10648_ (.CLK(clknet_leaf_103_clk),
    .D(_01279_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[31] ));
 sky130_fd_sc_hd__dfxtp_1 _10649_ (.CLK(clknet_leaf_79_clk),
    .D(_01280_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[32] ));
 sky130_fd_sc_hd__dfxtp_1 _10650_ (.CLK(clknet_leaf_80_clk),
    .D(_01281_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[33] ));
 sky130_fd_sc_hd__dfxtp_1 _10651_ (.CLK(clknet_leaf_80_clk),
    .D(_01282_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[34] ));
 sky130_fd_sc_hd__dfxtp_1 _10652_ (.CLK(clknet_leaf_79_clk),
    .D(_01283_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[35] ));
 sky130_fd_sc_hd__dfxtp_1 _10653_ (.CLK(clknet_leaf_80_clk),
    .D(_01284_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[36] ));
 sky130_fd_sc_hd__dfxtp_1 _10654_ (.CLK(clknet_leaf_81_clk),
    .D(_01285_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[37] ));
 sky130_fd_sc_hd__dfxtp_1 _10655_ (.CLK(clknet_leaf_81_clk),
    .D(_01286_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[38] ));
 sky130_fd_sc_hd__dfxtp_1 _10656_ (.CLK(clknet_leaf_82_clk),
    .D(_01287_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[39] ));
 sky130_fd_sc_hd__dfxtp_1 _10657_ (.CLK(clknet_leaf_66_clk),
    .D(_01288_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[40] ));
 sky130_fd_sc_hd__dfxtp_1 _10658_ (.CLK(clknet_leaf_67_clk),
    .D(_01289_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[41] ));
 sky130_fd_sc_hd__dfxtp_1 _10659_ (.CLK(clknet_leaf_67_clk),
    .D(_01290_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[42] ));
 sky130_fd_sc_hd__dfxtp_1 _10660_ (.CLK(clknet_leaf_67_clk),
    .D(_01291_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[43] ));
 sky130_fd_sc_hd__dfxtp_1 _10661_ (.CLK(clknet_leaf_66_clk),
    .D(_01292_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[44] ));
 sky130_fd_sc_hd__dfxtp_1 _10662_ (.CLK(clknet_leaf_68_clk),
    .D(_01293_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[45] ));
 sky130_fd_sc_hd__dfrtp_1 _10663_ (.CLK(clknet_leaf_106_clk),
    .D(_01294_),
    .RESET_B(_00053_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[96] ));
 sky130_fd_sc_hd__dfrtp_1 _10664_ (.CLK(clknet_leaf_106_clk),
    .D(_01295_),
    .RESET_B(_00054_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[97] ));
 sky130_fd_sc_hd__dfrtp_1 _10665_ (.CLK(clknet_leaf_106_clk),
    .D(_01296_),
    .RESET_B(_00055_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[98] ));
 sky130_fd_sc_hd__dfrtp_1 _10666_ (.CLK(clknet_leaf_106_clk),
    .D(_01297_),
    .RESET_B(_00056_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[99] ));
 sky130_fd_sc_hd__dfrtp_1 _10667_ (.CLK(clknet_leaf_110_clk),
    .D(_01298_),
    .RESET_B(_00057_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[100] ));
 sky130_fd_sc_hd__dfrtp_1 _10668_ (.CLK(clknet_leaf_110_clk),
    .D(_01299_),
    .RESET_B(_00058_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[101] ));
 sky130_fd_sc_hd__dfrtp_1 _10669_ (.CLK(clknet_leaf_98_clk),
    .D(_01300_),
    .RESET_B(_00059_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[102] ));
 sky130_fd_sc_hd__dfrtp_1 _10670_ (.CLK(clknet_leaf_110_clk),
    .D(_01301_),
    .RESET_B(_00060_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[103] ));
 sky130_fd_sc_hd__dfrtp_1 _10671_ (.CLK(clknet_leaf_106_clk),
    .D(_01302_),
    .RESET_B(_00061_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[104] ));
 sky130_fd_sc_hd__dfrtp_1 _10672_ (.CLK(clknet_leaf_106_clk),
    .D(_01303_),
    .RESET_B(_00062_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[105] ));
 sky130_fd_sc_hd__dfrtp_1 _10673_ (.CLK(clknet_leaf_106_clk),
    .D(_01304_),
    .RESET_B(_00063_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[106] ));
 sky130_fd_sc_hd__dfrtp_1 _10674_ (.CLK(clknet_leaf_110_clk),
    .D(_01305_),
    .RESET_B(_00064_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[107] ));
 sky130_fd_sc_hd__dfrtp_1 _10675_ (.CLK(clknet_leaf_109_clk),
    .D(_01306_),
    .RESET_B(_00065_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[108] ));
 sky130_fd_sc_hd__dfrtp_1 _10676_ (.CLK(clknet_leaf_107_clk),
    .D(_01307_),
    .RESET_B(_00066_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[109] ));
 sky130_fd_sc_hd__dfrtp_1 _10677_ (.CLK(clknet_leaf_108_clk),
    .D(_01308_),
    .RESET_B(_00067_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[110] ));
 sky130_fd_sc_hd__dfrtp_1 _10678_ (.CLK(clknet_leaf_108_clk),
    .D(_01309_),
    .RESET_B(_00068_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[111] ));
 sky130_fd_sc_hd__dfrtp_1 _10679_ (.CLK(clknet_leaf_11_clk),
    .D(_01310_),
    .RESET_B(_00069_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[112] ));
 sky130_fd_sc_hd__dfrtp_1 _10680_ (.CLK(clknet_leaf_116_clk),
    .D(_01311_),
    .RESET_B(_00070_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[113] ));
 sky130_fd_sc_hd__dfrtp_1 _10681_ (.CLK(clknet_leaf_3_clk),
    .D(_01312_),
    .RESET_B(_00071_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[114] ));
 sky130_fd_sc_hd__dfrtp_1 _10682_ (.CLK(clknet_leaf_3_clk),
    .D(_01313_),
    .RESET_B(_00072_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[115] ));
 sky130_fd_sc_hd__dfrtp_1 _10683_ (.CLK(clknet_leaf_116_clk),
    .D(_01314_),
    .RESET_B(_00073_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[116] ));
 sky130_fd_sc_hd__dfrtp_1 _10684_ (.CLK(clknet_leaf_3_clk),
    .D(_01315_),
    .RESET_B(_00074_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[117] ));
 sky130_fd_sc_hd__dfrtp_1 _10685_ (.CLK(clknet_leaf_108_clk),
    .D(_01316_),
    .RESET_B(_00075_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[118] ));
 sky130_fd_sc_hd__dfrtp_1 _10686_ (.CLK(clknet_leaf_108_clk),
    .D(_01317_),
    .RESET_B(_00076_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[119] ));
 sky130_fd_sc_hd__dfrtp_1 _10687_ (.CLK(clknet_leaf_11_clk),
    .D(_01318_),
    .RESET_B(_00077_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[120] ));
 sky130_fd_sc_hd__dfrtp_1 _10688_ (.CLK(clknet_leaf_11_clk),
    .D(_01319_),
    .RESET_B(_00078_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[121] ));
 sky130_fd_sc_hd__dfrtp_1 _10689_ (.CLK(clknet_leaf_107_clk),
    .D(_01320_),
    .RESET_B(_00079_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[122] ));
 sky130_fd_sc_hd__dfrtp_1 _10690_ (.CLK(clknet_leaf_107_clk),
    .D(_01321_),
    .RESET_B(_00080_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[123] ));
 sky130_fd_sc_hd__dfrtp_1 _10691_ (.CLK(clknet_leaf_108_clk),
    .D(_01322_),
    .RESET_B(_00081_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[124] ));
 sky130_fd_sc_hd__dfrtp_1 _10692_ (.CLK(clknet_leaf_108_clk),
    .D(_01323_),
    .RESET_B(_00082_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[125] ));
 sky130_fd_sc_hd__dfrtp_1 _10693_ (.CLK(clknet_leaf_107_clk),
    .D(_01324_),
    .RESET_B(_00083_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[126] ));
 sky130_fd_sc_hd__dfrtp_1 _10694_ (.CLK(clknet_leaf_107_clk),
    .D(_01325_),
    .RESET_B(_00084_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[127] ));
 sky130_fd_sc_hd__dfrtp_2 _10695_ (.CLK(clknet_leaf_21_clk),
    .D(_01326_),
    .RESET_B(_00085_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hist_addr[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10696_ (.CLK(clknet_leaf_21_clk),
    .D(_01327_),
    .RESET_B(_00086_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hist_addr[1] ));
 sky130_fd_sc_hd__dfrtp_1 _10697_ (.CLK(clknet_leaf_6_clk),
    .D(_01328_),
    .RESET_B(_00087_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hist_addr[2] ));
 sky130_fd_sc_hd__dfrtp_1 _10698_ (.CLK(clknet_leaf_7_clk),
    .D(net1613),
    .RESET_B(_00088_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hist_addr[3] ));
 sky130_fd_sc_hd__dfrtp_1 _10699_ (.CLK(clknet_leaf_21_clk),
    .D(_01330_),
    .RESET_B(_00089_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hist_addr[4] ));
 sky130_fd_sc_hd__dfrtp_1 _10700_ (.CLK(clknet_leaf_7_clk),
    .D(_01331_),
    .RESET_B(_00090_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hist_addr[5] ));
 sky130_fd_sc_hd__dfrtp_1 _10701_ (.CLK(clknet_leaf_7_clk),
    .D(_01332_),
    .RESET_B(_00091_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hist_addr[6] ));
 sky130_fd_sc_hd__dfrtp_1 _10702_ (.CLK(clknet_leaf_47_clk),
    .D(_01333_),
    .RESET_B(_00092_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.nulls[46] ));
 sky130_fd_sc_hd__dfrtp_1 _10703_ (.CLK(clknet_leaf_46_clk),
    .D(_01334_),
    .RESET_B(_00093_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.nulls[47] ));
 sky130_fd_sc_hd__dfrtp_1 _10704_ (.CLK(clknet_leaf_45_clk),
    .D(_01335_),
    .RESET_B(_00094_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.nulls[48] ));
 sky130_fd_sc_hd__dfrtp_1 _10705_ (.CLK(clknet_leaf_73_clk),
    .D(_01336_),
    .RESET_B(_00095_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.nulls[49] ));
 sky130_fd_sc_hd__dfrtp_1 _10706_ (.CLK(clknet_leaf_47_clk),
    .D(_01337_),
    .RESET_B(_00096_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.nulls[50] ));
 sky130_fd_sc_hd__dfrtp_1 _10707_ (.CLK(clknet_leaf_47_clk),
    .D(_01338_),
    .RESET_B(_00097_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.nulls[51] ));
 sky130_fd_sc_hd__dfrtp_1 _10708_ (.CLK(clknet_leaf_47_clk),
    .D(_01339_),
    .RESET_B(_00098_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.nulls[52] ));
 sky130_fd_sc_hd__dfrtp_1 _10709_ (.CLK(clknet_leaf_74_clk),
    .D(_01340_),
    .RESET_B(_00099_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.nulls[53] ));
 sky130_fd_sc_hd__dfrtp_1 _10710_ (.CLK(clknet_leaf_104_clk),
    .D(_01341_),
    .RESET_B(_00100_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.nulls[54] ));
 sky130_fd_sc_hd__dfrtp_1 _10711_ (.CLK(clknet_leaf_74_clk),
    .D(_01342_),
    .RESET_B(_00101_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.nulls[55] ));
 sky130_fd_sc_hd__dfrtp_1 _10712_ (.CLK(clknet_leaf_46_clk),
    .D(_01343_),
    .RESET_B(_00102_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.nulls[56] ));
 sky130_fd_sc_hd__dfrtp_1 _10713_ (.CLK(clknet_leaf_45_clk),
    .D(_01344_),
    .RESET_B(_00103_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.nulls[57] ));
 sky130_fd_sc_hd__dfrtp_1 _10714_ (.CLK(clknet_leaf_75_clk),
    .D(_01345_),
    .RESET_B(_00104_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.nulls[58] ));
 sky130_fd_sc_hd__dfrtp_1 _10715_ (.CLK(clknet_leaf_75_clk),
    .D(_01346_),
    .RESET_B(_00105_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.nulls[59] ));
 sky130_fd_sc_hd__dfrtp_1 _10716_ (.CLK(clknet_leaf_42_clk),
    .D(_01347_),
    .RESET_B(_00106_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.nulls[60] ));
 sky130_fd_sc_hd__dfrtp_1 _10717_ (.CLK(clknet_leaf_41_clk),
    .D(_01348_),
    .RESET_B(_00107_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.nulls[61] ));
 sky130_fd_sc_hd__dfrtp_1 _10718_ (.CLK(clknet_leaf_41_clk),
    .D(_01349_),
    .RESET_B(_00108_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.nulls[62] ));
 sky130_fd_sc_hd__dfrtp_1 _10719_ (.CLK(clknet_leaf_104_clk),
    .D(_01350_),
    .RESET_B(_00109_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.nulls[63] ));
 sky130_fd_sc_hd__dfrtp_1 _10720_ (.CLK(clknet_leaf_17_clk),
    .D(_01351_),
    .RESET_B(_00110_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.h_element[46] ));
 sky130_fd_sc_hd__dfrtp_1 _10721_ (.CLK(clknet_leaf_40_clk),
    .D(_01352_),
    .RESET_B(_00111_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.h_element[47] ));
 sky130_fd_sc_hd__dfrtp_1 _10722_ (.CLK(clknet_leaf_17_clk),
    .D(_01353_),
    .RESET_B(_00112_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.h_element[48] ));
 sky130_fd_sc_hd__dfrtp_1 _10723_ (.CLK(clknet_leaf_17_clk),
    .D(_01354_),
    .RESET_B(_00113_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.h_element[49] ));
 sky130_fd_sc_hd__dfrtp_1 _10724_ (.CLK(clknet_leaf_17_clk),
    .D(_01355_),
    .RESET_B(_00114_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.h_element[50] ));
 sky130_fd_sc_hd__dfrtp_1 _10725_ (.CLK(clknet_leaf_25_clk),
    .D(_01356_),
    .RESET_B(_00115_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.h_element[51] ));
 sky130_fd_sc_hd__dfrtp_1 _10726_ (.CLK(clknet_leaf_17_clk),
    .D(_01357_),
    .RESET_B(_00116_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.h_element[52] ));
 sky130_fd_sc_hd__dfrtp_1 _10727_ (.CLK(clknet_leaf_25_clk),
    .D(_01358_),
    .RESET_B(_00117_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.h_element[53] ));
 sky130_fd_sc_hd__dfrtp_2 _10728_ (.CLK(clknet_leaf_40_clk),
    .D(_01359_),
    .RESET_B(_00118_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.h_element[54] ));
 sky130_fd_sc_hd__dfrtp_1 _10729_ (.CLK(clknet_leaf_17_clk),
    .D(_01360_),
    .RESET_B(_00119_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.h_element[55] ));
 sky130_fd_sc_hd__dfrtp_1 _10730_ (.CLK(clknet_leaf_17_clk),
    .D(_01361_),
    .RESET_B(_00120_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.h_element[56] ));
 sky130_fd_sc_hd__dfrtp_1 _10731_ (.CLK(clknet_leaf_17_clk),
    .D(_01362_),
    .RESET_B(_00121_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.h_element[57] ));
 sky130_fd_sc_hd__dfrtp_1 _10732_ (.CLK(clknet_leaf_25_clk),
    .D(_01363_),
    .RESET_B(_00122_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.h_element[58] ));
 sky130_fd_sc_hd__dfrtp_1 _10733_ (.CLK(clknet_leaf_17_clk),
    .D(_01364_),
    .RESET_B(_00123_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.h_element[59] ));
 sky130_fd_sc_hd__dfrtp_1 _10734_ (.CLK(clknet_leaf_40_clk),
    .D(_01365_),
    .RESET_B(_00124_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.h_element[60] ));
 sky130_fd_sc_hd__dfrtp_1 _10735_ (.CLK(clknet_leaf_40_clk),
    .D(_01366_),
    .RESET_B(_00125_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.h_element[61] ));
 sky130_fd_sc_hd__dfrtp_1 _10736_ (.CLK(clknet_leaf_40_clk),
    .D(_01367_),
    .RESET_B(_00126_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.h_element[62] ));
 sky130_fd_sc_hd__dfrtp_1 _10737_ (.CLK(clknet_leaf_40_clk),
    .D(_01368_),
    .RESET_B(_00127_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.h_element[63] ));
 sky130_fd_sc_hd__dfstp_1 _10738_ (.CLK(clknet_leaf_5_clk),
    .D(_00028_),
    .SET_B(_00128_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10739_ (.CLK(clknet_leaf_4_clk),
    .D(_00029_),
    .RESET_B(_00129_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _10740_ (.CLK(clknet_leaf_4_clk),
    .D(_00030_),
    .RESET_B(_00130_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.state[2] ));
 sky130_fd_sc_hd__dfrtp_1 _10741_ (.CLK(clknet_leaf_6_clk),
    .D(_00031_),
    .RESET_B(_00131_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.state[3] ));
 sky130_fd_sc_hd__dfrtp_4 _10742_ (.CLK(clknet_leaf_6_clk),
    .D(_00032_),
    .RESET_B(_00132_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.eof_n ));
 sky130_fd_sc_hd__dfrtp_1 _10743_ (.CLK(clknet_leaf_6_clk),
    .D(_00033_),
    .RESET_B(_00133_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.state[5] ));
 sky130_fd_sc_hd__dfrtp_1 _10744_ (.CLK(clknet_leaf_6_clk),
    .D(_00034_),
    .RESET_B(_00134_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.state[6] ));
 sky130_fd_sc_hd__dfrtp_1 _10745_ (.CLK(clknet_leaf_6_clk),
    .D(net1480),
    .RESET_B(_00135_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.state[7] ));
 sky130_fd_sc_hd__dfstp_1 _10746_ (.CLK(clknet_leaf_6_clk),
    .D(_00036_),
    .SET_B(_00136_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.wr_r_en[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10747_ (.CLK(clknet_leaf_7_clk),
    .D(_00037_),
    .RESET_B(_00137_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.wr_r_en[1] ));
 sky130_fd_sc_hd__dfstp_2 _10748_ (.CLK(clknet_leaf_13_clk),
    .D(_00038_),
    .SET_B(_00138_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.sram_interface.word_cnt[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10749_ (.CLK(clknet_leaf_10_clk),
    .D(_00044_),
    .RESET_B(_00139_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.sram_interface.word_cnt[1] ));
 sky130_fd_sc_hd__dfrtp_4 _10750_ (.CLK(clknet_leaf_13_clk),
    .D(_00045_),
    .RESET_B(_00140_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.sram_interface.word_cnt[2] ));
 sky130_fd_sc_hd__dfrtp_4 _10751_ (.CLK(clknet_leaf_9_clk),
    .D(_00046_),
    .RESET_B(_00141_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.sram_interface.word_cnt[3] ));
 sky130_fd_sc_hd__dfrtp_1 _10752_ (.CLK(clknet_leaf_8_clk),
    .D(_00047_),
    .RESET_B(_00142_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.sram_interface.word_cnt[4] ));
 sky130_fd_sc_hd__dfrtp_1 _10753_ (.CLK(clknet_leaf_12_clk),
    .D(_00048_),
    .RESET_B(_00143_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.sram_interface.word_cnt[5] ));
 sky130_fd_sc_hd__dfrtp_1 _10754_ (.CLK(clknet_leaf_8_clk),
    .D(_00049_),
    .RESET_B(_00144_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.sram_interface.word_cnt[6] ));
 sky130_fd_sc_hd__dfrtp_1 _10755_ (.CLK(clknet_leaf_10_clk),
    .D(_00050_),
    .RESET_B(_00145_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.sram_interface.word_cnt[7] ));
 sky130_fd_sc_hd__dfrtp_1 _10756_ (.CLK(clknet_leaf_10_clk),
    .D(_00051_),
    .RESET_B(_00146_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.sram_interface.word_cnt[8] ));
 sky130_fd_sc_hd__dfrtp_2 _10757_ (.CLK(clknet_leaf_13_clk),
    .D(_00052_),
    .RESET_B(_00147_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.sram_interface.word_cnt[9] ));
 sky130_fd_sc_hd__dfrtp_1 _10758_ (.CLK(clknet_leaf_12_clk),
    .D(_00039_),
    .RESET_B(_00148_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.sram_interface.word_cnt[10] ));
 sky130_fd_sc_hd__dfrtp_1 _10759_ (.CLK(clknet_leaf_8_clk),
    .D(net1041),
    .RESET_B(_00149_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.sram_interface.word_cnt[11] ));
 sky130_fd_sc_hd__dfrtp_1 _10760_ (.CLK(clknet_leaf_9_clk),
    .D(_00041_),
    .RESET_B(_00150_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.sram_interface.word_cnt[12] ));
 sky130_fd_sc_hd__dfrtp_2 _10761_ (.CLK(clknet_leaf_9_clk),
    .D(_00042_),
    .RESET_B(_00151_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.sram_interface.word_cnt[13] ));
 sky130_fd_sc_hd__dfrtp_1 _10762_ (.CLK(clknet_leaf_12_clk),
    .D(_00043_),
    .RESET_B(_00152_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.sram_interface.word_cnt[14] ));
 sky130_fd_sc_hd__dfrtp_1 _10763_ (.CLK(clknet_leaf_111_clk),
    .D(_01369_),
    .RESET_B(_00153_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[64] ));
 sky130_fd_sc_hd__dfrtp_1 _10764_ (.CLK(clknet_leaf_111_clk),
    .D(_01370_),
    .RESET_B(_00154_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[65] ));
 sky130_fd_sc_hd__dfrtp_1 _10765_ (.CLK(clknet_leaf_97_clk),
    .D(_01371_),
    .RESET_B(_00155_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[66] ));
 sky130_fd_sc_hd__dfrtp_1 _10766_ (.CLK(clknet_leaf_111_clk),
    .D(_01372_),
    .RESET_B(_00156_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[67] ));
 sky130_fd_sc_hd__dfrtp_1 _10767_ (.CLK(clknet_leaf_110_clk),
    .D(_01373_),
    .RESET_B(_00157_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[68] ));
 sky130_fd_sc_hd__dfrtp_1 _10768_ (.CLK(clknet_leaf_111_clk),
    .D(_01374_),
    .RESET_B(_00158_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[69] ));
 sky130_fd_sc_hd__dfrtp_1 _10769_ (.CLK(clknet_leaf_111_clk),
    .D(_01375_),
    .RESET_B(_00159_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[70] ));
 sky130_fd_sc_hd__dfrtp_1 _10770_ (.CLK(clknet_leaf_111_clk),
    .D(_01376_),
    .RESET_B(_00160_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[71] ));
 sky130_fd_sc_hd__dfrtp_1 _10771_ (.CLK(clknet_leaf_111_clk),
    .D(_01377_),
    .RESET_B(_00161_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[72] ));
 sky130_fd_sc_hd__dfrtp_1 _10772_ (.CLK(clknet_leaf_113_clk),
    .D(_01378_),
    .RESET_B(_00162_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[73] ));
 sky130_fd_sc_hd__dfrtp_1 _10773_ (.CLK(clknet_leaf_113_clk),
    .D(_01379_),
    .RESET_B(_00163_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[74] ));
 sky130_fd_sc_hd__dfrtp_1 _10774_ (.CLK(clknet_leaf_113_clk),
    .D(_01380_),
    .RESET_B(_00164_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[75] ));
 sky130_fd_sc_hd__dfrtp_1 _10775_ (.CLK(clknet_leaf_109_clk),
    .D(_01381_),
    .RESET_B(_00165_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[76] ));
 sky130_fd_sc_hd__dfrtp_1 _10776_ (.CLK(clknet_leaf_109_clk),
    .D(_01382_),
    .RESET_B(_00166_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[77] ));
 sky130_fd_sc_hd__dfrtp_1 _10777_ (.CLK(clknet_leaf_113_clk),
    .D(_01383_),
    .RESET_B(_00167_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[78] ));
 sky130_fd_sc_hd__dfrtp_1 _10778_ (.CLK(clknet_leaf_113_clk),
    .D(_01384_),
    .RESET_B(_00168_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[79] ));
 sky130_fd_sc_hd__dfrtp_1 _10779_ (.CLK(clknet_leaf_118_clk),
    .D(_01385_),
    .RESET_B(_00169_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[80] ));
 sky130_fd_sc_hd__dfrtp_1 _10780_ (.CLK(clknet_leaf_118_clk),
    .D(_01386_),
    .RESET_B(_00170_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[81] ));
 sky130_fd_sc_hd__dfrtp_1 _10781_ (.CLK(clknet_leaf_118_clk),
    .D(_01387_),
    .RESET_B(_00171_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[82] ));
 sky130_fd_sc_hd__dfrtp_1 _10782_ (.CLK(clknet_leaf_118_clk),
    .D(_01388_),
    .RESET_B(_00172_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[83] ));
 sky130_fd_sc_hd__dfrtp_1 _10783_ (.CLK(clknet_leaf_117_clk),
    .D(_01389_),
    .RESET_B(_00173_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[84] ));
 sky130_fd_sc_hd__dfrtp_1 _10784_ (.CLK(clknet_leaf_117_clk),
    .D(_01390_),
    .RESET_B(_00174_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[85] ));
 sky130_fd_sc_hd__dfrtp_1 _10785_ (.CLK(clknet_leaf_114_clk),
    .D(_01391_),
    .RESET_B(_00175_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[86] ));
 sky130_fd_sc_hd__dfrtp_1 _10786_ (.CLK(clknet_leaf_114_clk),
    .D(_01392_),
    .RESET_B(_00176_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[87] ));
 sky130_fd_sc_hd__dfrtp_1 _10787_ (.CLK(clknet_leaf_117_clk),
    .D(_01393_),
    .RESET_B(_00177_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[88] ));
 sky130_fd_sc_hd__dfrtp_1 _10788_ (.CLK(clknet_leaf_117_clk),
    .D(_01394_),
    .RESET_B(_00178_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[89] ));
 sky130_fd_sc_hd__dfrtp_1 _10789_ (.CLK(clknet_leaf_117_clk),
    .D(_01395_),
    .RESET_B(_00179_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[90] ));
 sky130_fd_sc_hd__dfrtp_1 _10790_ (.CLK(clknet_leaf_117_clk),
    .D(_01396_),
    .RESET_B(_00180_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[91] ));
 sky130_fd_sc_hd__dfrtp_1 _10791_ (.CLK(clknet_leaf_114_clk),
    .D(_01397_),
    .RESET_B(_00181_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[92] ));
 sky130_fd_sc_hd__dfrtp_1 _10792_ (.CLK(clknet_leaf_114_clk),
    .D(_01398_),
    .RESET_B(_00182_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[93] ));
 sky130_fd_sc_hd__dfrtp_1 _10793_ (.CLK(clknet_leaf_113_clk),
    .D(_01399_),
    .RESET_B(_00183_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[94] ));
 sky130_fd_sc_hd__dfrtp_1 _10794_ (.CLK(clknet_leaf_113_clk),
    .D(_01400_),
    .RESET_B(_00184_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[95] ));
 sky130_fd_sc_hd__dfstp_1 _10795_ (.CLK(clknet_leaf_4_clk),
    .D(_00000_),
    .SET_B(_00185_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.WB.curr_state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10796_ (.CLK(clknet_leaf_3_clk),
    .D(_00001_),
    .RESET_B(_00186_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.WB.curr_state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _10797_ (.CLK(clknet_leaf_3_clk),
    .D(_00002_),
    .RESET_B(_00187_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.WB.curr_state[2] ));
 sky130_fd_sc_hd__dfrtp_4 _10798_ (.CLK(clknet_leaf_18_clk),
    .D(_01401_),
    .RESET_B(_00188_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.max_index[1] ));
 sky130_fd_sc_hd__dfrtp_4 _10799_ (.CLK(clknet_leaf_18_clk),
    .D(_01402_),
    .RESET_B(_00189_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.max_index[2] ));
 sky130_fd_sc_hd__dfrtp_2 _10800_ (.CLK(clknet_leaf_17_clk),
    .D(_01403_),
    .RESET_B(_00190_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.max_index[3] ));
 sky130_fd_sc_hd__dfrtp_2 _10801_ (.CLK(clknet_leaf_18_clk),
    .D(_01404_),
    .RESET_B(_00191_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.max_index[4] ));
 sky130_fd_sc_hd__dfrtp_4 _10802_ (.CLK(clknet_leaf_20_clk),
    .D(_01405_),
    .RESET_B(_00192_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.max_index[5] ));
 sky130_fd_sc_hd__dfrtp_2 _10803_ (.CLK(clknet_leaf_18_clk),
    .D(_01406_),
    .RESET_B(_00193_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.max_index[6] ));
 sky130_fd_sc_hd__dfrtp_2 _10804_ (.CLK(clknet_leaf_18_clk),
    .D(_01407_),
    .RESET_B(_00194_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.max_index[7] ));
 sky130_fd_sc_hd__dfstp_1 _10805_ (.CLK(clknet_leaf_25_clk),
    .D(_00003_),
    .SET_B(_00195_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.curr_state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10806_ (.CLK(clknet_leaf_39_clk),
    .D(_00004_),
    .RESET_B(_00196_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.curr_state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _10807_ (.CLK(clknet_leaf_31_clk),
    .D(_00005_),
    .RESET_B(_00197_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.curr_state[2] ));
 sky130_fd_sc_hd__dfrtp_1 _10808_ (.CLK(clknet_leaf_26_clk),
    .D(_00006_),
    .RESET_B(_00198_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.finished ));
 sky130_fd_sc_hd__dfrtp_1 _10809_ (.CLK(clknet_leaf_32_clk),
    .D(_00007_),
    .RESET_B(_00199_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.curr_state[4] ));
 sky130_fd_sc_hd__dfrtp_1 _10810_ (.CLK(clknet_leaf_39_clk),
    .D(_00008_),
    .RESET_B(_00200_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.curr_state[5] ));
 sky130_fd_sc_hd__dfrtp_4 _10811_ (.CLK(clknet_leaf_32_clk),
    .D(_00009_),
    .RESET_B(_00201_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10812_ (.CLK(clknet_leaf_26_clk),
    .D(_00010_),
    .RESET_B(_00202_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.pulse_first_n ));
 sky130_fd_sc_hd__dfrtp_1 _10813_ (.CLK(clknet_leaf_25_clk),
    .D(_00011_),
    .RESET_B(_00203_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.curr_state[8] ));
 sky130_fd_sc_hd__dfrtp_1 _10814_ (.CLK(clknet_leaf_111_clk),
    .D(_01408_),
    .RESET_B(_00204_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10815_ (.CLK(clknet_leaf_111_clk),
    .D(_01409_),
    .RESET_B(_00205_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[1] ));
 sky130_fd_sc_hd__dfrtp_1 _10816_ (.CLK(clknet_leaf_97_clk),
    .D(_01410_),
    .RESET_B(_00206_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[2] ));
 sky130_fd_sc_hd__dfrtp_1 _10817_ (.CLK(clknet_leaf_98_clk),
    .D(_01411_),
    .RESET_B(_00207_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[3] ));
 sky130_fd_sc_hd__dfrtp_1 _10818_ (.CLK(clknet_leaf_97_clk),
    .D(_01412_),
    .RESET_B(_00208_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[4] ));
 sky130_fd_sc_hd__dfrtp_1 _10819_ (.CLK(clknet_leaf_97_clk),
    .D(_01413_),
    .RESET_B(_00209_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[5] ));
 sky130_fd_sc_hd__dfrtp_1 _10820_ (.CLK(clknet_leaf_97_clk),
    .D(_01414_),
    .RESET_B(_00210_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[6] ));
 sky130_fd_sc_hd__dfrtp_1 _10821_ (.CLK(clknet_leaf_97_clk),
    .D(_01415_),
    .RESET_B(_00211_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[7] ));
 sky130_fd_sc_hd__dfrtp_1 _10822_ (.CLK(clknet_leaf_111_clk),
    .D(_01416_),
    .RESET_B(_00212_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[8] ));
 sky130_fd_sc_hd__dfrtp_1 _10823_ (.CLK(clknet_leaf_97_clk),
    .D(_01417_),
    .RESET_B(_00213_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[9] ));
 sky130_fd_sc_hd__dfrtp_1 _10824_ (.CLK(clknet_leaf_97_clk),
    .D(_01418_),
    .RESET_B(_00214_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[10] ));
 sky130_fd_sc_hd__dfrtp_1 _10825_ (.CLK(clknet_leaf_97_clk),
    .D(_01419_),
    .RESET_B(_00215_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[11] ));
 sky130_fd_sc_hd__dfrtp_1 _10826_ (.CLK(clknet_leaf_112_clk),
    .D(_01420_),
    .RESET_B(_00216_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[12] ));
 sky130_fd_sc_hd__dfrtp_1 _10827_ (.CLK(clknet_leaf_113_clk),
    .D(_01421_),
    .RESET_B(_00217_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[13] ));
 sky130_fd_sc_hd__dfrtp_1 _10828_ (.CLK(clknet_leaf_96_clk),
    .D(_01422_),
    .RESET_B(_00218_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[14] ));
 sky130_fd_sc_hd__dfrtp_1 _10829_ (.CLK(clknet_leaf_97_clk),
    .D(_01423_),
    .RESET_B(_00219_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[15] ));
 sky130_fd_sc_hd__dfrtp_1 _10830_ (.CLK(clknet_leaf_116_clk),
    .D(_01424_),
    .RESET_B(_00220_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[16] ));
 sky130_fd_sc_hd__dfrtp_1 _10831_ (.CLK(clknet_leaf_116_clk),
    .D(_01425_),
    .RESET_B(_00221_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[17] ));
 sky130_fd_sc_hd__dfrtp_1 _10832_ (.CLK(clknet_leaf_117_clk),
    .D(_01426_),
    .RESET_B(_00222_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[18] ));
 sky130_fd_sc_hd__dfrtp_1 _10833_ (.CLK(clknet_leaf_117_clk),
    .D(_01427_),
    .RESET_B(_00223_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[19] ));
 sky130_fd_sc_hd__dfrtp_1 _10834_ (.CLK(clknet_leaf_116_clk),
    .D(_01428_),
    .RESET_B(_00224_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[20] ));
 sky130_fd_sc_hd__dfrtp_1 _10835_ (.CLK(clknet_leaf_116_clk),
    .D(_01429_),
    .RESET_B(_00225_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[21] ));
 sky130_fd_sc_hd__dfrtp_1 _10836_ (.CLK(clknet_leaf_115_clk),
    .D(_01430_),
    .RESET_B(_00226_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[22] ));
 sky130_fd_sc_hd__dfrtp_1 _10837_ (.CLK(clknet_leaf_115_clk),
    .D(_01431_),
    .RESET_B(_00227_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[23] ));
 sky130_fd_sc_hd__dfrtp_1 _10838_ (.CLK(clknet_leaf_115_clk),
    .D(_01432_),
    .RESET_B(_00228_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[24] ));
 sky130_fd_sc_hd__dfrtp_1 _10839_ (.CLK(clknet_leaf_116_clk),
    .D(_01433_),
    .RESET_B(_00229_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[25] ));
 sky130_fd_sc_hd__dfrtp_1 _10840_ (.CLK(clknet_leaf_116_clk),
    .D(_01434_),
    .RESET_B(_00230_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[26] ));
 sky130_fd_sc_hd__dfrtp_1 _10841_ (.CLK(clknet_leaf_116_clk),
    .D(_01435_),
    .RESET_B(_00231_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[27] ));
 sky130_fd_sc_hd__dfrtp_1 _10842_ (.CLK(clknet_leaf_108_clk),
    .D(_01436_),
    .RESET_B(_00232_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[28] ));
 sky130_fd_sc_hd__dfrtp_1 _10843_ (.CLK(clknet_leaf_108_clk),
    .D(_01437_),
    .RESET_B(_00233_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[29] ));
 sky130_fd_sc_hd__dfrtp_1 _10844_ (.CLK(clknet_leaf_108_clk),
    .D(_01438_),
    .RESET_B(_00234_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[30] ));
 sky130_fd_sc_hd__dfrtp_1 _10845_ (.CLK(clknet_leaf_108_clk),
    .D(_01439_),
    .RESET_B(_00235_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[31] ));
 sky130_fd_sc_hd__dfstp_1 _10846_ (.CLK(clknet_leaf_2_clk),
    .D(_01440_),
    .SET_B(_00236_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.translation.totalEn ));
 sky130_fd_sc_hd__dfrtp_1 _10847_ (.CLK(clknet_leaf_2_clk),
    .D(_01441_),
    .RESET_B(_00237_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.translation.resEn ));
 sky130_fd_sc_hd__dfstp_1 _10848_ (.CLK(clknet_leaf_117_clk),
    .D(_01442_),
    .SET_B(_00238_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.translation.index[0] ));
 sky130_fd_sc_hd__dfstp_1 _10849_ (.CLK(clknet_leaf_117_clk),
    .D(_01443_),
    .SET_B(_00239_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.translation.index[1] ));
 sky130_fd_sc_hd__dfstp_1 _10850_ (.CLK(clknet_leaf_2_clk),
    .D(_01444_),
    .SET_B(_00240_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.translation.index[2] ));
 sky130_fd_sc_hd__dfstp_1 _10851_ (.CLK(clknet_leaf_2_clk),
    .D(_01445_),
    .SET_B(_00241_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.translation.index[3] ));
 sky130_fd_sc_hd__dfstp_1 _10852_ (.CLK(clknet_leaf_116_clk),
    .D(_01446_),
    .SET_B(_00242_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.translation.index[4] ));
 sky130_fd_sc_hd__dfrtp_4 _10853_ (.CLK(clknet_leaf_116_clk),
    .D(_01447_),
    .RESET_B(_00243_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.translation.index[5] ));
 sky130_fd_sc_hd__dfrtp_4 _10854_ (.CLK(clknet_leaf_116_clk),
    .D(_01448_),
    .RESET_B(_00244_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.translation.index[6] ));
 sky130_fd_sc_hd__dfrtp_1 _10855_ (.CLK(clknet_leaf_2_clk),
    .D(_01449_),
    .RESET_B(_00245_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.translation.writeEn ));
 sky130_fd_sc_hd__dfrtp_1 _10856_ (.CLK(clknet_leaf_11_clk),
    .D(_01450_),
    .RESET_B(_00246_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.sram_interface.TRN_counter[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10857_ (.CLK(clknet_leaf_11_clk),
    .D(_01451_),
    .RESET_B(_00247_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.sram_interface.TRN_counter[1] ));
 sky130_fd_sc_hd__dfrtp_1 _10858_ (.CLK(clknet_leaf_10_clk),
    .D(_01452_),
    .RESET_B(_00248_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.sram_interface.TRN_counter[2] ));
 sky130_fd_sc_hd__dfrtp_1 _10859_ (.CLK(clknet_leaf_28_clk),
    .D(\top.header_synthesis.next_zero_count[0] ),
    .RESET_B(_00249_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.zero_count[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10860_ (.CLK(clknet_leaf_28_clk),
    .D(\top.header_synthesis.next_zero_count[1] ),
    .RESET_B(_00250_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.zero_count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _10861_ (.CLK(clknet_leaf_29_clk),
    .D(\top.header_synthesis.next_zero_count[2] ),
    .RESET_B(_00251_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.zero_count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _10862_ (.CLK(clknet_leaf_29_clk),
    .D(\top.header_synthesis.next_zero_count[3] ),
    .RESET_B(_00252_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.zero_count[3] ));
 sky130_fd_sc_hd__dfrtp_1 _10863_ (.CLK(clknet_leaf_28_clk),
    .D(\top.header_synthesis.next_zero_count[4] ),
    .RESET_B(_00253_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.zero_count[4] ));
 sky130_fd_sc_hd__dfrtp_1 _10864_ (.CLK(clknet_leaf_28_clk),
    .D(\top.header_synthesis.next_zero_count[5] ),
    .RESET_B(_00254_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.zero_count[5] ));
 sky130_fd_sc_hd__dfrtp_1 _10865_ (.CLK(clknet_leaf_28_clk),
    .D(\top.header_synthesis.next_zero_count[6] ),
    .RESET_B(_00255_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.zero_count[6] ));
 sky130_fd_sc_hd__dfrtp_1 _10866_ (.CLK(clknet_leaf_28_clk),
    .D(\top.header_synthesis.next_zero_count[7] ),
    .RESET_B(_00256_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.zero_count[7] ));
 sky130_fd_sc_hd__dfstp_1 _10867_ (.CLK(clknet_leaf_14_clk),
    .D(_01453_),
    .SET_B(_00257_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.finish_check ));
 sky130_fd_sc_hd__dfrtp_4 _10868_ (.CLK(clknet_leaf_26_clk),
    .D(\top.header_synthesis.next_enable ),
    .RESET_B(_00258_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.header_synthesis.enable ));
 sky130_fd_sc_hd__dfrtp_1 _10869_ (.CLK(clknet_leaf_27_clk),
    .D(_01454_),
    .RESET_B(_00259_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.header_synthesis.count[0] ));
 sky130_fd_sc_hd__dfrtp_2 _10870_ (.CLK(clknet_leaf_27_clk),
    .D(_01455_),
    .RESET_B(_00260_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.header_synthesis.count[1] ));
 sky130_fd_sc_hd__dfrtp_2 _10871_ (.CLK(clknet_leaf_27_clk),
    .D(_01456_),
    .RESET_B(_00261_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.header_synthesis.count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _10872_ (.CLK(clknet_leaf_27_clk),
    .D(_01457_),
    .RESET_B(_00262_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.header_synthesis.count[3] ));
 sky130_fd_sc_hd__dfrtp_1 _10873_ (.CLK(clknet_leaf_27_clk),
    .D(_01458_),
    .RESET_B(_00263_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.header_synthesis.count[4] ));
 sky130_fd_sc_hd__dfrtp_1 _10874_ (.CLK(clknet_leaf_23_clk),
    .D(_01459_),
    .RESET_B(_00264_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.header_synthesis.count[5] ));
 sky130_fd_sc_hd__dfrtp_1 _10875_ (.CLK(clknet_leaf_23_clk),
    .D(_01460_),
    .RESET_B(_00265_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.header_synthesis.count[6] ));
 sky130_fd_sc_hd__dfrtp_1 _10876_ (.CLK(clknet_leaf_23_clk),
    .D(_01461_),
    .RESET_B(_00266_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.header_synthesis.count[7] ));
 sky130_fd_sc_hd__dfrtp_1 _10877_ (.CLK(clknet_leaf_26_clk),
    .D(\top.header_synthesis.next_char_added ),
    .RESET_B(_00267_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.header_synthesis.char_added ));
 sky130_fd_sc_hd__dfrtp_1 _10878_ (.CLK(clknet_leaf_23_clk),
    .D(\top.header_synthesis.next_header[0] ),
    .RESET_B(_00268_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.header_synthesis.header[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10879_ (.CLK(clknet_leaf_24_clk),
    .D(\top.header_synthesis.next_header[1] ),
    .RESET_B(_00269_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.header_synthesis.header[1] ));
 sky130_fd_sc_hd__dfrtp_1 _10880_ (.CLK(clknet_leaf_23_clk),
    .D(\top.header_synthesis.next_header[2] ),
    .RESET_B(_00270_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.header_synthesis.header[2] ));
 sky130_fd_sc_hd__dfrtp_1 _10881_ (.CLK(clknet_leaf_23_clk),
    .D(\top.header_synthesis.next_header[3] ),
    .RESET_B(_00271_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.header_synthesis.header[3] ));
 sky130_fd_sc_hd__dfrtp_1 _10882_ (.CLK(clknet_leaf_23_clk),
    .D(\top.header_synthesis.next_header[4] ),
    .RESET_B(_00272_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.header_synthesis.header[4] ));
 sky130_fd_sc_hd__dfrtp_1 _10883_ (.CLK(clknet_leaf_23_clk),
    .D(\top.header_synthesis.next_header[5] ),
    .RESET_B(_00273_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.header_synthesis.header[5] ));
 sky130_fd_sc_hd__dfrtp_1 _10884_ (.CLK(clknet_leaf_23_clk),
    .D(\top.header_synthesis.next_header[6] ),
    .RESET_B(_00274_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.header_synthesis.header[6] ));
 sky130_fd_sc_hd__dfrtp_1 _10885_ (.CLK(clknet_leaf_23_clk),
    .D(\top.header_synthesis.next_header[7] ),
    .RESET_B(_00275_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.header_synthesis.header[7] ));
 sky130_fd_sc_hd__dfrtp_1 _10886_ (.CLK(clknet_leaf_23_clk),
    .D(\top.header_synthesis.next_header[8] ),
    .RESET_B(_00276_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.header_synthesis.header[8] ));
 sky130_fd_sc_hd__dfrtp_1 _10887_ (.CLK(clknet_leaf_26_clk),
    .D(\top.header_synthesis.next_start ),
    .RESET_B(_00277_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.header_synthesis.start ));
 sky130_fd_sc_hd__dfrtp_1 _10888_ (.CLK(clknet_leaf_28_clk),
    .D(\top.header_synthesis.next_write_zeroes ),
    .RESET_B(_00278_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.header_synthesis.write_zeroes ));
 sky130_fd_sc_hd__dfrtp_1 _10889_ (.CLK(clknet_leaf_26_clk),
    .D(\top.header_synthesis.next_write_char_path ),
    .RESET_B(_00279_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.header_synthesis.write_char_path ));
 sky130_fd_sc_hd__dfrtp_1 _10890_ (.CLK(clknet_leaf_32_clk),
    .D(_01462_),
    .RESET_B(_00280_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.pulse_first ));
 sky130_fd_sc_hd__dfrtp_1 _10891_ (.CLK(clknet_leaf_33_clk),
    .D(net1483),
    .RESET_B(_00281_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.end_cond ));
 sky130_fd_sc_hd__dfrtp_4 _10892_ (.CLK(clknet_leaf_31_clk),
    .D(_01464_),
    .RESET_B(_00282_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.i[0] ));
 sky130_fd_sc_hd__dfrtp_2 _10893_ (.CLK(clknet_leaf_31_clk),
    .D(_01465_),
    .RESET_B(_00283_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.i[1] ));
 sky130_fd_sc_hd__dfrtp_2 _10894_ (.CLK(clknet_leaf_34_clk),
    .D(_01466_),
    .RESET_B(_00284_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.i[2] ));
 sky130_fd_sc_hd__dfrtp_1 _10895_ (.CLK(clknet_leaf_31_clk),
    .D(_01467_),
    .RESET_B(_00285_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.i[3] ));
 sky130_fd_sc_hd__dfrtp_1 _10896_ (.CLK(clknet_leaf_31_clk),
    .D(_01468_),
    .RESET_B(_00286_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.i[4] ));
 sky130_fd_sc_hd__dfrtp_1 _10897_ (.CLK(clknet_leaf_31_clk),
    .D(_01469_),
    .RESET_B(_00287_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.i[5] ));
 sky130_fd_sc_hd__dfrtp_1 _10898_ (.CLK(clknet_leaf_33_clk),
    .D(_01470_),
    .RESET_B(_00288_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.i[6] ));
 sky130_fd_sc_hd__dfrtp_1 _10899_ (.CLK(clknet_leaf_33_clk),
    .D(_01471_),
    .RESET_B(_00289_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.cb_enable ));
 sky130_fd_sc_hd__dfstp_1 _10900_ (.CLK(clknet_leaf_51_clk),
    .D(_01472_),
    .SET_B(_00290_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.end_cnt[0] ));
 sky130_fd_sc_hd__dfstp_1 _10901_ (.CLK(clknet_leaf_51_clk),
    .D(_01473_),
    .SET_B(_00291_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.end_cnt[1] ));
 sky130_fd_sc_hd__dfstp_1 _10902_ (.CLK(clknet_leaf_50_clk),
    .D(_01474_),
    .SET_B(_00292_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.end_cnt[2] ));
 sky130_fd_sc_hd__dfstp_2 _10903_ (.CLK(clknet_leaf_51_clk),
    .D(_01475_),
    .SET_B(_00293_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.end_cnt[3] ));
 sky130_fd_sc_hd__dfstp_2 _10904_ (.CLK(clknet_leaf_51_clk),
    .D(_01476_),
    .SET_B(_00294_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.end_cnt[4] ));
 sky130_fd_sc_hd__dfstp_1 _10905_ (.CLK(clknet_leaf_37_clk),
    .D(_01477_),
    .SET_B(_00295_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.end_cnt[5] ));
 sky130_fd_sc_hd__dfstp_1 _10906_ (.CLK(clknet_leaf_33_clk),
    .D(_01478_),
    .SET_B(_00296_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.end_cnt[6] ));
 sky130_fd_sc_hd__dfrtp_1 _10907_ (.CLK(clknet_leaf_32_clk),
    .D(_01479_),
    .RESET_B(_00297_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.check_right ));
 sky130_fd_sc_hd__dfrtp_1 _10908_ (.CLK(clknet_leaf_33_clk),
    .D(_01480_),
    .RESET_B(_00298_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.end_check ));
 sky130_fd_sc_hd__dfrtp_1 _10909_ (.CLK(clknet_leaf_3_clk),
    .D(\top.controller.fin_TRN ),
    .RESET_B(_00299_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.controller.fin_reg[1] ));
 sky130_fd_sc_hd__dfrtp_2 _10910_ (.CLK(clknet_leaf_25_clk),
    .D(net954),
    .RESET_B(_00300_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.controller.fin_reg[2] ));
 sky130_fd_sc_hd__dfrtp_1 _10911_ (.CLK(clknet_leaf_11_clk),
    .D(net977),
    .RESET_B(_00301_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.controller.fin_reg[3] ));
 sky130_fd_sc_hd__dfrtp_1 _10912_ (.CLK(clknet_leaf_106_clk),
    .D(net953),
    .RESET_B(_00302_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.controller.fin_reg[4] ));
 sky130_fd_sc_hd__dfrtp_1 _10913_ (.CLK(clknet_leaf_107_clk),
    .D(net955),
    .RESET_B(_00303_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.controller.fin_reg[5] ));
 sky130_fd_sc_hd__dfrtp_1 _10914_ (.CLK(clknet_leaf_4_clk),
    .D(net952),
    .RESET_B(_00304_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.controller.fin_reg[6] ));
 sky130_fd_sc_hd__dfrtp_1 _10915_ (.CLK(clknet_leaf_5_clk),
    .D(net918),
    .RESET_B(_00305_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.controller.fin_reg[7] ));
 sky130_fd_sc_hd__dfrtp_1 _10916_ (.CLK(clknet_leaf_33_clk),
    .D(_01481_),
    .RESET_B(_00306_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.left_check ));
 sky130_fd_sc_hd__dfrtp_1 _10917_ (.CLK(clknet_leaf_39_clk),
    .D(_01482_),
    .RESET_B(_00307_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_found ));
 sky130_fd_sc_hd__dfrtp_1 _10918_ (.CLK(clknet_leaf_46_clk),
    .D(_01483_),
    .RESET_B(_00308_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10919_ (.CLK(clknet_leaf_48_clk),
    .D(_01484_),
    .RESET_B(_00309_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[1] ));
 sky130_fd_sc_hd__dfrtp_1 _10920_ (.CLK(clknet_leaf_47_clk),
    .D(_01485_),
    .RESET_B(_00310_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[2] ));
 sky130_fd_sc_hd__dfrtp_1 _10921_ (.CLK(clknet_leaf_71_clk),
    .D(_01486_),
    .RESET_B(_00311_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[3] ));
 sky130_fd_sc_hd__dfrtp_1 _10922_ (.CLK(clknet_leaf_71_clk),
    .D(_01487_),
    .RESET_B(_00312_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[4] ));
 sky130_fd_sc_hd__dfrtp_1 _10923_ (.CLK(clknet_leaf_71_clk),
    .D(_01488_),
    .RESET_B(_00313_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[5] ));
 sky130_fd_sc_hd__dfrtp_1 _10924_ (.CLK(clknet_leaf_71_clk),
    .D(_01489_),
    .RESET_B(_00314_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[6] ));
 sky130_fd_sc_hd__dfrtp_1 _10925_ (.CLK(clknet_leaf_65_clk),
    .D(_01490_),
    .RESET_B(_00315_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[7] ));
 sky130_fd_sc_hd__dfrtp_1 _10926_ (.CLK(clknet_leaf_61_clk),
    .D(_01491_),
    .RESET_B(_00316_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[8] ));
 sky130_fd_sc_hd__dfrtp_1 _10927_ (.CLK(clknet_leaf_61_clk),
    .D(_01492_),
    .RESET_B(_00317_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[9] ));
 sky130_fd_sc_hd__dfrtp_1 _10928_ (.CLK(clknet_leaf_61_clk),
    .D(_01493_),
    .RESET_B(_00318_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[10] ));
 sky130_fd_sc_hd__dfrtp_1 _10929_ (.CLK(clknet_leaf_60_clk),
    .D(_01494_),
    .RESET_B(_00319_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[11] ));
 sky130_fd_sc_hd__dfrtp_1 _10930_ (.CLK(clknet_leaf_60_clk),
    .D(_01495_),
    .RESET_B(_00320_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[12] ));
 sky130_fd_sc_hd__dfrtp_1 _10931_ (.CLK(clknet_leaf_59_clk),
    .D(_01496_),
    .RESET_B(_00321_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[13] ));
 sky130_fd_sc_hd__dfrtp_1 _10932_ (.CLK(clknet_leaf_59_clk),
    .D(_01497_),
    .RESET_B(_00322_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[14] ));
 sky130_fd_sc_hd__dfrtp_1 _10933_ (.CLK(clknet_leaf_58_clk),
    .D(_01498_),
    .RESET_B(_00323_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[15] ));
 sky130_fd_sc_hd__dfrtp_1 _10934_ (.CLK(clknet_leaf_58_clk),
    .D(_01499_),
    .RESET_B(_00324_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[16] ));
 sky130_fd_sc_hd__dfrtp_1 _10935_ (.CLK(clknet_leaf_58_clk),
    .D(net1199),
    .RESET_B(_00325_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[17] ));
 sky130_fd_sc_hd__dfrtp_1 _10936_ (.CLK(clknet_leaf_54_clk),
    .D(_01501_),
    .RESET_B(_00326_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[18] ));
 sky130_fd_sc_hd__dfrtp_1 _10937_ (.CLK(clknet_leaf_54_clk),
    .D(_01502_),
    .RESET_B(_00327_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[19] ));
 sky130_fd_sc_hd__dfrtp_1 _10938_ (.CLK(clknet_leaf_55_clk),
    .D(_01503_),
    .RESET_B(_00328_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[20] ));
 sky130_fd_sc_hd__dfrtp_1 _10939_ (.CLK(clknet_leaf_53_clk),
    .D(_01504_),
    .RESET_B(_00329_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[21] ));
 sky130_fd_sc_hd__dfrtp_1 _10940_ (.CLK(clknet_leaf_52_clk),
    .D(_01505_),
    .RESET_B(_00330_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[22] ));
 sky130_fd_sc_hd__dfrtp_1 _10941_ (.CLK(clknet_leaf_51_clk),
    .D(_01506_),
    .RESET_B(_00331_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[23] ));
 sky130_fd_sc_hd__dfrtp_1 _10942_ (.CLK(clknet_leaf_52_clk),
    .D(_01507_),
    .RESET_B(_00332_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[24] ));
 sky130_fd_sc_hd__dfrtp_1 _10943_ (.CLK(clknet_leaf_37_clk),
    .D(_01508_),
    .RESET_B(_00333_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[25] ));
 sky130_fd_sc_hd__dfrtp_1 _10944_ (.CLK(clknet_leaf_36_clk),
    .D(_01509_),
    .RESET_B(_00334_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[26] ));
 sky130_fd_sc_hd__dfrtp_1 _10945_ (.CLK(clknet_leaf_37_clk),
    .D(_01510_),
    .RESET_B(_00335_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[27] ));
 sky130_fd_sc_hd__dfrtp_1 _10946_ (.CLK(clknet_leaf_35_clk),
    .D(_01511_),
    .RESET_B(_00336_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[28] ));
 sky130_fd_sc_hd__dfrtp_1 _10947_ (.CLK(clknet_leaf_38_clk),
    .D(net1427),
    .RESET_B(_00337_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[29] ));
 sky130_fd_sc_hd__dfrtp_1 _10948_ (.CLK(clknet_leaf_39_clk),
    .D(_01513_),
    .RESET_B(_00338_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[30] ));
 sky130_fd_sc_hd__dfrtp_1 _10949_ (.CLK(clknet_leaf_41_clk),
    .D(_01514_),
    .RESET_B(_00339_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[31] ));
 sky130_fd_sc_hd__dfrtp_1 _10950_ (.CLK(clknet_leaf_46_clk),
    .D(_01515_),
    .RESET_B(_00340_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[32] ));
 sky130_fd_sc_hd__dfrtp_1 _10951_ (.CLK(clknet_leaf_47_clk),
    .D(_01516_),
    .RESET_B(_00341_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[33] ));
 sky130_fd_sc_hd__dfrtp_1 _10952_ (.CLK(clknet_leaf_47_clk),
    .D(net1355),
    .RESET_B(_00342_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[34] ));
 sky130_fd_sc_hd__dfrtp_1 _10953_ (.CLK(clknet_leaf_70_clk),
    .D(_01518_),
    .RESET_B(_00343_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[35] ));
 sky130_fd_sc_hd__dfrtp_1 _10954_ (.CLK(clknet_leaf_70_clk),
    .D(_01519_),
    .RESET_B(_00344_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[36] ));
 sky130_fd_sc_hd__dfrtp_1 _10955_ (.CLK(clknet_leaf_64_clk),
    .D(_01520_),
    .RESET_B(_00345_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[37] ));
 sky130_fd_sc_hd__dfrtp_1 _10956_ (.CLK(clknet_leaf_64_clk),
    .D(_01521_),
    .RESET_B(_00346_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[38] ));
 sky130_fd_sc_hd__dfrtp_1 _10957_ (.CLK(clknet_leaf_65_clk),
    .D(_01522_),
    .RESET_B(_00347_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[39] ));
 sky130_fd_sc_hd__dfrtp_1 _10958_ (.CLK(clknet_leaf_65_clk),
    .D(_01523_),
    .RESET_B(_00348_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[40] ));
 sky130_fd_sc_hd__dfrtp_1 _10959_ (.CLK(clknet_leaf_62_clk),
    .D(_01524_),
    .RESET_B(_00349_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[41] ));
 sky130_fd_sc_hd__dfrtp_1 _10960_ (.CLK(clknet_leaf_61_clk),
    .D(net1361),
    .RESET_B(_00350_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[42] ));
 sky130_fd_sc_hd__dfrtp_1 _10961_ (.CLK(clknet_leaf_61_clk),
    .D(_01526_),
    .RESET_B(_00351_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[43] ));
 sky130_fd_sc_hd__dfrtp_1 _10962_ (.CLK(clknet_leaf_61_clk),
    .D(_01527_),
    .RESET_B(_00352_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[44] ));
 sky130_fd_sc_hd__dfrtp_1 _10963_ (.CLK(clknet_leaf_61_clk),
    .D(_01528_),
    .RESET_B(_00353_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[45] ));
 sky130_fd_sc_hd__dfrtp_1 _10964_ (.CLK(clknet_leaf_57_clk),
    .D(_01529_),
    .RESET_B(_00354_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[46] ));
 sky130_fd_sc_hd__dfrtp_1 _10965_ (.CLK(clknet_leaf_56_clk),
    .D(_01530_),
    .RESET_B(_00355_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[47] ));
 sky130_fd_sc_hd__dfrtp_1 _10966_ (.CLK(clknet_leaf_56_clk),
    .D(_01531_),
    .RESET_B(_00356_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[48] ));
 sky130_fd_sc_hd__dfrtp_1 _10967_ (.CLK(clknet_leaf_56_clk),
    .D(_01532_),
    .RESET_B(_00357_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[49] ));
 sky130_fd_sc_hd__dfrtp_1 _10968_ (.CLK(clknet_leaf_55_clk),
    .D(net1130),
    .RESET_B(_00358_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[50] ));
 sky130_fd_sc_hd__dfrtp_1 _10969_ (.CLK(clknet_leaf_55_clk),
    .D(net1122),
    .RESET_B(_00359_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[51] ));
 sky130_fd_sc_hd__dfrtp_1 _10970_ (.CLK(clknet_leaf_55_clk),
    .D(net1137),
    .RESET_B(_00360_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[52] ));
 sky130_fd_sc_hd__dfrtp_1 _10971_ (.CLK(clknet_leaf_48_clk),
    .D(net1072),
    .RESET_B(_00361_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[53] ));
 sky130_fd_sc_hd__dfrtp_1 _10972_ (.CLK(clknet_leaf_48_clk),
    .D(_01537_),
    .RESET_B(_00362_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[54] ));
 sky130_fd_sc_hd__dfrtp_1 _10973_ (.CLK(clknet_leaf_49_clk),
    .D(_01538_),
    .RESET_B(_00363_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[55] ));
 sky130_fd_sc_hd__dfrtp_1 _10974_ (.CLK(clknet_leaf_50_clk),
    .D(_01539_),
    .RESET_B(_00364_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[56] ));
 sky130_fd_sc_hd__dfrtp_1 _10975_ (.CLK(clknet_leaf_37_clk),
    .D(_01540_),
    .RESET_B(_00365_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[57] ));
 sky130_fd_sc_hd__dfrtp_1 _10976_ (.CLK(clknet_leaf_37_clk),
    .D(_01541_),
    .RESET_B(_00366_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[58] ));
 sky130_fd_sc_hd__dfrtp_1 _10977_ (.CLK(clknet_leaf_37_clk),
    .D(_01542_),
    .RESET_B(_00367_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[59] ));
 sky130_fd_sc_hd__dfrtp_1 _10978_ (.CLK(clknet_leaf_38_clk),
    .D(_01543_),
    .RESET_B(_00368_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[60] ));
 sky130_fd_sc_hd__dfrtp_1 _10979_ (.CLK(clknet_leaf_38_clk),
    .D(_01544_),
    .RESET_B(_00369_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[61] ));
 sky130_fd_sc_hd__dfrtp_1 _10980_ (.CLK(clknet_leaf_39_clk),
    .D(_01545_),
    .RESET_B(_00370_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[62] ));
 sky130_fd_sc_hd__dfrtp_1 _10981_ (.CLK(clknet_leaf_39_clk),
    .D(_01546_),
    .RESET_B(_00371_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[63] ));
 sky130_fd_sc_hd__dfrtp_1 _10982_ (.CLK(clknet_leaf_42_clk),
    .D(_01547_),
    .RESET_B(_00372_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[64] ));
 sky130_fd_sc_hd__dfrtp_1 _10983_ (.CLK(clknet_leaf_47_clk),
    .D(net1386),
    .RESET_B(_00373_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[65] ));
 sky130_fd_sc_hd__dfrtp_1 _10984_ (.CLK(clknet_leaf_47_clk),
    .D(net1424),
    .RESET_B(_00374_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[66] ));
 sky130_fd_sc_hd__dfrtp_1 _10985_ (.CLK(clknet_leaf_71_clk),
    .D(_01550_),
    .RESET_B(_00375_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[67] ));
 sky130_fd_sc_hd__dfrtp_1 _10986_ (.CLK(clknet_leaf_71_clk),
    .D(_01551_),
    .RESET_B(_00376_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[68] ));
 sky130_fd_sc_hd__dfrtp_1 _10987_ (.CLK(clknet_leaf_70_clk),
    .D(_01552_),
    .RESET_B(_00377_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[69] ));
 sky130_fd_sc_hd__dfrtp_1 _10988_ (.CLK(clknet_leaf_70_clk),
    .D(net1178),
    .RESET_B(_00378_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[70] ));
 sky130_fd_sc_hd__dfrtp_1 _10989_ (.CLK(clknet_leaf_65_clk),
    .D(net1348),
    .RESET_B(_00379_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[71] ));
 sky130_fd_sc_hd__dfrtp_1 _10990_ (.CLK(clknet_leaf_65_clk),
    .D(_01555_),
    .RESET_B(_00380_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[72] ));
 sky130_fd_sc_hd__dfrtp_1 _10991_ (.CLK(clknet_leaf_62_clk),
    .D(_01556_),
    .RESET_B(_00381_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[73] ));
 sky130_fd_sc_hd__dfrtp_1 _10992_ (.CLK(clknet_leaf_61_clk),
    .D(_01557_),
    .RESET_B(_00382_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[74] ));
 sky130_fd_sc_hd__dfrtp_1 _10993_ (.CLK(clknet_leaf_60_clk),
    .D(_01558_),
    .RESET_B(_00383_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[75] ));
 sky130_fd_sc_hd__dfrtp_1 _10994_ (.CLK(clknet_leaf_60_clk),
    .D(net1540),
    .RESET_B(_00384_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[76] ));
 sky130_fd_sc_hd__dfrtp_1 _10995_ (.CLK(clknet_leaf_59_clk),
    .D(_01560_),
    .RESET_B(_00385_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[77] ));
 sky130_fd_sc_hd__dfrtp_1 _10996_ (.CLK(clknet_leaf_58_clk),
    .D(_01561_),
    .RESET_B(_00386_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[78] ));
 sky130_fd_sc_hd__dfrtp_1 _10997_ (.CLK(clknet_leaf_58_clk),
    .D(_01562_),
    .RESET_B(_00387_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[79] ));
 sky130_fd_sc_hd__dfrtp_1 _10998_ (.CLK(clknet_leaf_58_clk),
    .D(net1113),
    .RESET_B(_00388_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[80] ));
 sky130_fd_sc_hd__dfrtp_1 _10999_ (.CLK(clknet_leaf_54_clk),
    .D(net1246),
    .RESET_B(_00389_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[81] ));
 sky130_fd_sc_hd__dfrtp_1 _11000_ (.CLK(clknet_leaf_54_clk),
    .D(_01565_),
    .RESET_B(_00390_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[82] ));
 sky130_fd_sc_hd__dfrtp_1 _11001_ (.CLK(clknet_leaf_53_clk),
    .D(_01566_),
    .RESET_B(_00391_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[83] ));
 sky130_fd_sc_hd__dfrtp_1 _11002_ (.CLK(clknet_leaf_54_clk),
    .D(_01567_),
    .RESET_B(_00392_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[84] ));
 sky130_fd_sc_hd__dfrtp_1 _11003_ (.CLK(clknet_leaf_53_clk),
    .D(_01568_),
    .RESET_B(_00393_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[85] ));
 sky130_fd_sc_hd__dfrtp_1 _11004_ (.CLK(clknet_leaf_52_clk),
    .D(_01569_),
    .RESET_B(_00394_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[86] ));
 sky130_fd_sc_hd__dfrtp_1 _11005_ (.CLK(clknet_leaf_52_clk),
    .D(_01570_),
    .RESET_B(_00395_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[87] ));
 sky130_fd_sc_hd__dfrtp_1 _11006_ (.CLK(clknet_leaf_52_clk),
    .D(_01571_),
    .RESET_B(_00396_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[88] ));
 sky130_fd_sc_hd__dfrtp_1 _11007_ (.CLK(clknet_leaf_36_clk),
    .D(_01572_),
    .RESET_B(_00397_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[89] ));
 sky130_fd_sc_hd__dfrtp_1 _11008_ (.CLK(clknet_leaf_36_clk),
    .D(_01573_),
    .RESET_B(_00398_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[90] ));
 sky130_fd_sc_hd__dfrtp_1 _11009_ (.CLK(clknet_leaf_35_clk),
    .D(net1440),
    .RESET_B(_00399_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[91] ));
 sky130_fd_sc_hd__dfrtp_1 _11010_ (.CLK(clknet_leaf_35_clk),
    .D(_01575_),
    .RESET_B(_00400_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[92] ));
 sky130_fd_sc_hd__dfrtp_1 _11011_ (.CLK(clknet_leaf_38_clk),
    .D(net1293),
    .RESET_B(_00401_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[93] ));
 sky130_fd_sc_hd__dfrtp_1 _11012_ (.CLK(clknet_leaf_39_clk),
    .D(_01577_),
    .RESET_B(_00402_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[94] ));
 sky130_fd_sc_hd__dfrtp_1 _11013_ (.CLK(clknet_leaf_41_clk),
    .D(net1330),
    .RESET_B(_00403_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[95] ));
 sky130_fd_sc_hd__dfrtp_1 _11014_ (.CLK(clknet_leaf_46_clk),
    .D(_01579_),
    .RESET_B(_00404_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[96] ));
 sky130_fd_sc_hd__dfrtp_1 _11015_ (.CLK(clknet_leaf_47_clk),
    .D(_01580_),
    .RESET_B(_00405_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[97] ));
 sky130_fd_sc_hd__dfrtp_1 _11016_ (.CLK(clknet_leaf_47_clk),
    .D(_01581_),
    .RESET_B(_00406_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[98] ));
 sky130_fd_sc_hd__dfrtp_1 _11017_ (.CLK(clknet_leaf_63_clk),
    .D(_01582_),
    .RESET_B(_00407_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[99] ));
 sky130_fd_sc_hd__dfrtp_1 _11018_ (.CLK(clknet_leaf_70_clk),
    .D(net1214),
    .RESET_B(_00408_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[100] ));
 sky130_fd_sc_hd__dfrtp_1 _11019_ (.CLK(clknet_leaf_64_clk),
    .D(_01584_),
    .RESET_B(_00409_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[101] ));
 sky130_fd_sc_hd__dfrtp_1 _11020_ (.CLK(clknet_leaf_64_clk),
    .D(_01585_),
    .RESET_B(_00410_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[102] ));
 sky130_fd_sc_hd__dfrtp_1 _11021_ (.CLK(clknet_leaf_64_clk),
    .D(_01586_),
    .RESET_B(_00411_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[103] ));
 sky130_fd_sc_hd__dfrtp_1 _11022_ (.CLK(clknet_leaf_65_clk),
    .D(_01587_),
    .RESET_B(_00412_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[104] ));
 sky130_fd_sc_hd__dfrtp_1 _11023_ (.CLK(clknet_leaf_62_clk),
    .D(_01588_),
    .RESET_B(_00413_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[105] ));
 sky130_fd_sc_hd__dfrtp_1 _11024_ (.CLK(clknet_leaf_61_clk),
    .D(_01589_),
    .RESET_B(_00414_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[106] ));
 sky130_fd_sc_hd__dfrtp_1 _11025_ (.CLK(clknet_leaf_61_clk),
    .D(_01590_),
    .RESET_B(_00415_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[107] ));
 sky130_fd_sc_hd__dfrtp_1 _11026_ (.CLK(clknet_leaf_60_clk),
    .D(_01591_),
    .RESET_B(_00416_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[108] ));
 sky130_fd_sc_hd__dfrtp_1 _11027_ (.CLK(clknet_leaf_60_clk),
    .D(_01592_),
    .RESET_B(_00417_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[109] ));
 sky130_fd_sc_hd__dfrtp_1 _11028_ (.CLK(clknet_leaf_57_clk),
    .D(_01593_),
    .RESET_B(_00418_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[110] ));
 sky130_fd_sc_hd__dfrtp_1 _11029_ (.CLK(clknet_leaf_56_clk),
    .D(net1098),
    .RESET_B(_00419_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[111] ));
 sky130_fd_sc_hd__dfrtp_1 _11030_ (.CLK(clknet_leaf_57_clk),
    .D(_01595_),
    .RESET_B(_00420_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[112] ));
 sky130_fd_sc_hd__dfrtp_1 _11031_ (.CLK(clknet_leaf_55_clk),
    .D(_01596_),
    .RESET_B(_00421_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[113] ));
 sky130_fd_sc_hd__dfrtp_1 _11032_ (.CLK(clknet_leaf_55_clk),
    .D(_01597_),
    .RESET_B(_00422_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[114] ));
 sky130_fd_sc_hd__dfrtp_1 _11033_ (.CLK(clknet_leaf_55_clk),
    .D(_01598_),
    .RESET_B(_00423_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[115] ));
 sky130_fd_sc_hd__dfrtp_1 _11034_ (.CLK(clknet_leaf_55_clk),
    .D(_01599_),
    .RESET_B(_00424_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[116] ));
 sky130_fd_sc_hd__dfrtp_1 _11035_ (.CLK(clknet_leaf_49_clk),
    .D(net1273),
    .RESET_B(_00425_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[117] ));
 sky130_fd_sc_hd__dfrtp_1 _11036_ (.CLK(clknet_leaf_49_clk),
    .D(_01601_),
    .RESET_B(_00426_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[118] ));
 sky130_fd_sc_hd__dfrtp_1 _11037_ (.CLK(clknet_leaf_51_clk),
    .D(_01602_),
    .RESET_B(_00427_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[119] ));
 sky130_fd_sc_hd__dfrtp_1 _11038_ (.CLK(clknet_leaf_50_clk),
    .D(_01603_),
    .RESET_B(_00428_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[120] ));
 sky130_fd_sc_hd__dfrtp_1 _11039_ (.CLK(clknet_leaf_37_clk),
    .D(_01604_),
    .RESET_B(_00429_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[121] ));
 sky130_fd_sc_hd__dfrtp_1 _11040_ (.CLK(clknet_leaf_37_clk),
    .D(_01605_),
    .RESET_B(_00430_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[122] ));
 sky130_fd_sc_hd__dfrtp_1 _11041_ (.CLK(clknet_leaf_37_clk),
    .D(_01606_),
    .RESET_B(_00431_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[123] ));
 sky130_fd_sc_hd__dfrtp_1 _11042_ (.CLK(clknet_leaf_38_clk),
    .D(_01607_),
    .RESET_B(_00432_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[124] ));
 sky130_fd_sc_hd__dfrtp_1 _11043_ (.CLK(clknet_leaf_38_clk),
    .D(_01608_),
    .RESET_B(_00433_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[125] ));
 sky130_fd_sc_hd__dfrtp_1 _11044_ (.CLK(clknet_leaf_39_clk),
    .D(_01609_),
    .RESET_B(_00434_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[126] ));
 sky130_fd_sc_hd__dfrtp_1 _11045_ (.CLK(clknet_leaf_39_clk),
    .D(_01610_),
    .RESET_B(_00435_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path[127] ));
 sky130_fd_sc_hd__dfrtp_1 _11046_ (.CLK(clknet_leaf_24_clk),
    .D(_01611_),
    .RESET_B(_00436_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_index[0] ));
 sky130_fd_sc_hd__dfrtp_4 _11047_ (.CLK(clknet_leaf_24_clk),
    .D(_01612_),
    .RESET_B(_00437_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_index[1] ));
 sky130_fd_sc_hd__dfrtp_4 _11048_ (.CLK(clknet_leaf_24_clk),
    .D(_01613_),
    .RESET_B(_00438_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_index[2] ));
 sky130_fd_sc_hd__dfrtp_4 _11049_ (.CLK(clknet_leaf_24_clk),
    .D(_01614_),
    .RESET_B(_00439_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_index[3] ));
 sky130_fd_sc_hd__dfrtp_2 _11050_ (.CLK(clknet_leaf_24_clk),
    .D(_01615_),
    .RESET_B(_00440_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_index[4] ));
 sky130_fd_sc_hd__dfrtp_2 _11051_ (.CLK(clknet_leaf_24_clk),
    .D(_01616_),
    .RESET_B(_00441_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_index[5] ));
 sky130_fd_sc_hd__dfrtp_4 _11052_ (.CLK(clknet_leaf_24_clk),
    .D(_01617_),
    .RESET_B(_00442_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_index[6] ));
 sky130_fd_sc_hd__dfrtp_1 _11053_ (.CLK(clknet_leaf_25_clk),
    .D(_01618_),
    .RESET_B(_00443_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_index[7] ));
 sky130_fd_sc_hd__dfrtp_1 _11054_ (.CLK(clknet_leaf_32_clk),
    .D(_01619_),
    .RESET_B(_00444_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.state8 ));
 sky130_fd_sc_hd__dfstp_2 _11055_ (.CLK(clknet_leaf_39_clk),
    .D(_01620_),
    .SET_B(_00445_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[1] ));
 sky130_fd_sc_hd__dfrtp_4 _11056_ (.CLK(clknet_leaf_48_clk),
    .D(_01621_),
    .RESET_B(_00446_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11057_ (.CLK(clknet_leaf_48_clk),
    .D(_01622_),
    .RESET_B(_00447_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11058_ (.CLK(clknet_leaf_47_clk),
    .D(_01623_),
    .RESET_B(_00448_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[4] ));
 sky130_fd_sc_hd__dfrtp_1 _11059_ (.CLK(clknet_leaf_71_clk),
    .D(_01624_),
    .RESET_B(_00449_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[5] ));
 sky130_fd_sc_hd__dfrtp_2 _11060_ (.CLK(clknet_leaf_48_clk),
    .D(_01625_),
    .RESET_B(_00450_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[6] ));
 sky130_fd_sc_hd__dfrtp_2 _11061_ (.CLK(clknet_leaf_56_clk),
    .D(_01626_),
    .RESET_B(_00451_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[7] ));
 sky130_fd_sc_hd__dfrtp_2 _11062_ (.CLK(clknet_leaf_61_clk),
    .D(_01627_),
    .RESET_B(_00452_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[8] ));
 sky130_fd_sc_hd__dfrtp_2 _11063_ (.CLK(clknet_leaf_61_clk),
    .D(_01628_),
    .RESET_B(_00453_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[9] ));
 sky130_fd_sc_hd__dfrtp_2 _11064_ (.CLK(clknet_leaf_60_clk),
    .D(_01629_),
    .RESET_B(_00454_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[10] ));
 sky130_fd_sc_hd__dfrtp_2 _11065_ (.CLK(clknet_leaf_60_clk),
    .D(_01630_),
    .RESET_B(_00455_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[11] ));
 sky130_fd_sc_hd__dfrtp_1 _11066_ (.CLK(clknet_leaf_60_clk),
    .D(_01631_),
    .RESET_B(_00456_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[12] ));
 sky130_fd_sc_hd__dfrtp_1 _11067_ (.CLK(clknet_leaf_59_clk),
    .D(_01632_),
    .RESET_B(_00457_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[13] ));
 sky130_fd_sc_hd__dfrtp_1 _11068_ (.CLK(clknet_leaf_59_clk),
    .D(_01633_),
    .RESET_B(_00458_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[14] ));
 sky130_fd_sc_hd__dfrtp_1 _11069_ (.CLK(clknet_leaf_58_clk),
    .D(_01634_),
    .RESET_B(_00459_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[15] ));
 sky130_fd_sc_hd__dfrtp_1 _11070_ (.CLK(clknet_leaf_57_clk),
    .D(_01635_),
    .RESET_B(_00460_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[16] ));
 sky130_fd_sc_hd__dfrtp_2 _11071_ (.CLK(clknet_leaf_57_clk),
    .D(_01636_),
    .RESET_B(_00461_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[17] ));
 sky130_fd_sc_hd__dfrtp_1 _11072_ (.CLK(clknet_leaf_54_clk),
    .D(_01637_),
    .RESET_B(_00462_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[18] ));
 sky130_fd_sc_hd__dfrtp_1 _11073_ (.CLK(clknet_leaf_53_clk),
    .D(_01638_),
    .RESET_B(_00463_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[19] ));
 sky130_fd_sc_hd__dfrtp_1 _11074_ (.CLK(clknet_leaf_53_clk),
    .D(_01639_),
    .RESET_B(_00464_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[20] ));
 sky130_fd_sc_hd__dfrtp_1 _11075_ (.CLK(clknet_leaf_52_clk),
    .D(_01640_),
    .RESET_B(_00465_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[21] ));
 sky130_fd_sc_hd__dfrtp_2 _11076_ (.CLK(clknet_leaf_52_clk),
    .D(_01641_),
    .RESET_B(_00466_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[22] ));
 sky130_fd_sc_hd__dfrtp_2 _11077_ (.CLK(clknet_leaf_52_clk),
    .D(_01642_),
    .RESET_B(_00467_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[23] ));
 sky130_fd_sc_hd__dfrtp_2 _11078_ (.CLK(clknet_leaf_52_clk),
    .D(_01643_),
    .RESET_B(_00468_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[24] ));
 sky130_fd_sc_hd__dfrtp_2 _11079_ (.CLK(clknet_leaf_52_clk),
    .D(_01644_),
    .RESET_B(_00469_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[25] ));
 sky130_fd_sc_hd__dfrtp_1 _11080_ (.CLK(clknet_leaf_52_clk),
    .D(_01645_),
    .RESET_B(_00470_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[26] ));
 sky130_fd_sc_hd__dfrtp_1 _11081_ (.CLK(clknet_leaf_36_clk),
    .D(_01646_),
    .RESET_B(_00471_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[27] ));
 sky130_fd_sc_hd__dfrtp_1 _11082_ (.CLK(clknet_leaf_36_clk),
    .D(_01647_),
    .RESET_B(_00472_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[28] ));
 sky130_fd_sc_hd__dfrtp_2 _11083_ (.CLK(clknet_leaf_36_clk),
    .D(_01648_),
    .RESET_B(_00473_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[29] ));
 sky130_fd_sc_hd__dfrtp_2 _11084_ (.CLK(clknet_leaf_37_clk),
    .D(_01649_),
    .RESET_B(_00474_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[30] ));
 sky130_fd_sc_hd__dfrtp_2 _11085_ (.CLK(clknet_leaf_37_clk),
    .D(_01650_),
    .RESET_B(_00475_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[31] ));
 sky130_fd_sc_hd__dfrtp_2 _11086_ (.CLK(clknet_leaf_42_clk),
    .D(_01651_),
    .RESET_B(_00476_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[32] ));
 sky130_fd_sc_hd__dfrtp_4 _11087_ (.CLK(clknet_leaf_46_clk),
    .D(_01652_),
    .RESET_B(_00477_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[33] ));
 sky130_fd_sc_hd__dfrtp_2 _11088_ (.CLK(clknet_leaf_63_clk),
    .D(_01653_),
    .RESET_B(_00478_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[34] ));
 sky130_fd_sc_hd__dfrtp_1 _11089_ (.CLK(clknet_leaf_63_clk),
    .D(_01654_),
    .RESET_B(_00479_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[35] ));
 sky130_fd_sc_hd__dfrtp_1 _11090_ (.CLK(clknet_leaf_63_clk),
    .D(_01655_),
    .RESET_B(_00480_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[36] ));
 sky130_fd_sc_hd__dfrtp_2 _11091_ (.CLK(clknet_leaf_63_clk),
    .D(_01656_),
    .RESET_B(_00481_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[37] ));
 sky130_fd_sc_hd__dfrtp_2 _11092_ (.CLK(clknet_leaf_64_clk),
    .D(_01657_),
    .RESET_B(_00482_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[38] ));
 sky130_fd_sc_hd__dfrtp_2 _11093_ (.CLK(clknet_leaf_65_clk),
    .D(_01658_),
    .RESET_B(_00483_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[39] ));
 sky130_fd_sc_hd__dfrtp_2 _11094_ (.CLK(clknet_leaf_62_clk),
    .D(_01659_),
    .RESET_B(_00484_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[40] ));
 sky130_fd_sc_hd__dfrtp_1 _11095_ (.CLK(clknet_leaf_62_clk),
    .D(_01660_),
    .RESET_B(_00485_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[41] ));
 sky130_fd_sc_hd__dfrtp_2 _11096_ (.CLK(clknet_leaf_62_clk),
    .D(_01661_),
    .RESET_B(_00486_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[42] ));
 sky130_fd_sc_hd__dfrtp_2 _11097_ (.CLK(clknet_leaf_61_clk),
    .D(_01662_),
    .RESET_B(_00487_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[43] ));
 sky130_fd_sc_hd__dfrtp_2 _11098_ (.CLK(clknet_leaf_61_clk),
    .D(_01663_),
    .RESET_B(_00488_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[44] ));
 sky130_fd_sc_hd__dfrtp_1 _11099_ (.CLK(clknet_leaf_62_clk),
    .D(_01664_),
    .RESET_B(_00489_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[45] ));
 sky130_fd_sc_hd__dfrtp_1 _11100_ (.CLK(clknet_leaf_62_clk),
    .D(_01665_),
    .RESET_B(_00490_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[46] ));
 sky130_fd_sc_hd__dfrtp_1 _11101_ (.CLK(clknet_leaf_56_clk),
    .D(_01666_),
    .RESET_B(_00491_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[47] ));
 sky130_fd_sc_hd__dfrtp_1 _11102_ (.CLK(clknet_leaf_56_clk),
    .D(_01667_),
    .RESET_B(_00492_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[48] ));
 sky130_fd_sc_hd__dfrtp_2 _11103_ (.CLK(clknet_leaf_56_clk),
    .D(_01668_),
    .RESET_B(_00493_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[49] ));
 sky130_fd_sc_hd__dfrtp_2 _11104_ (.CLK(clknet_leaf_56_clk),
    .D(_01669_),
    .RESET_B(_00494_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[50] ));
 sky130_fd_sc_hd__dfrtp_2 _11105_ (.CLK(clknet_leaf_56_clk),
    .D(_01670_),
    .RESET_B(_00495_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[51] ));
 sky130_fd_sc_hd__dfrtp_2 _11106_ (.CLK(clknet_leaf_48_clk),
    .D(_01671_),
    .RESET_B(_00496_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[52] ));
 sky130_fd_sc_hd__dfrtp_2 _11107_ (.CLK(clknet_leaf_48_clk),
    .D(_01672_),
    .RESET_B(_00497_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[53] ));
 sky130_fd_sc_hd__dfrtp_1 _11108_ (.CLK(clknet_leaf_49_clk),
    .D(_01673_),
    .RESET_B(_00498_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[54] ));
 sky130_fd_sc_hd__dfrtp_1 _11109_ (.CLK(clknet_leaf_49_clk),
    .D(_01674_),
    .RESET_B(_00499_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[55] ));
 sky130_fd_sc_hd__dfrtp_1 _11110_ (.CLK(clknet_leaf_49_clk),
    .D(_01675_),
    .RESET_B(_00500_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[56] ));
 sky130_fd_sc_hd__dfrtp_1 _11111_ (.CLK(clknet_leaf_50_clk),
    .D(_01676_),
    .RESET_B(_00501_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[57] ));
 sky130_fd_sc_hd__dfrtp_1 _11112_ (.CLK(clknet_leaf_50_clk),
    .D(_01677_),
    .RESET_B(_00502_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[58] ));
 sky130_fd_sc_hd__dfrtp_2 _11113_ (.CLK(clknet_leaf_37_clk),
    .D(_01678_),
    .RESET_B(_00503_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[59] ));
 sky130_fd_sc_hd__dfrtp_1 _11114_ (.CLK(clknet_leaf_38_clk),
    .D(_01679_),
    .RESET_B(_00504_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[60] ));
 sky130_fd_sc_hd__dfrtp_1 _11115_ (.CLK(clknet_leaf_38_clk),
    .D(_01680_),
    .RESET_B(_00505_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[61] ));
 sky130_fd_sc_hd__dfrtp_2 _11116_ (.CLK(clknet_leaf_38_clk),
    .D(_01681_),
    .RESET_B(_00506_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[62] ));
 sky130_fd_sc_hd__dfrtp_2 _11117_ (.CLK(clknet_leaf_50_clk),
    .D(_01682_),
    .RESET_B(_00507_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[63] ));
 sky130_fd_sc_hd__dfrtp_1 _11118_ (.CLK(clknet_leaf_50_clk),
    .D(_01683_),
    .RESET_B(_00508_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[64] ));
 sky130_fd_sc_hd__dfrtp_2 _11119_ (.CLK(clknet_leaf_49_clk),
    .D(_01684_),
    .RESET_B(_00509_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[65] ));
 sky130_fd_sc_hd__dfrtp_2 _11120_ (.CLK(clknet_leaf_63_clk),
    .D(_01685_),
    .RESET_B(_00510_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[66] ));
 sky130_fd_sc_hd__dfrtp_1 _11121_ (.CLK(clknet_leaf_63_clk),
    .D(_01686_),
    .RESET_B(_00511_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[67] ));
 sky130_fd_sc_hd__dfrtp_1 _11122_ (.CLK(clknet_leaf_71_clk),
    .D(_01687_),
    .RESET_B(_00512_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[68] ));
 sky130_fd_sc_hd__dfrtp_2 _11123_ (.CLK(clknet_leaf_70_clk),
    .D(_01688_),
    .RESET_B(_00513_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[69] ));
 sky130_fd_sc_hd__dfrtp_2 _11124_ (.CLK(clknet_leaf_56_clk),
    .D(_01689_),
    .RESET_B(_00514_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[70] ));
 sky130_fd_sc_hd__dfrtp_2 _11125_ (.CLK(clknet_leaf_62_clk),
    .D(_01690_),
    .RESET_B(_00515_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[71] ));
 sky130_fd_sc_hd__dfrtp_2 _11126_ (.CLK(clknet_leaf_61_clk),
    .D(_01691_),
    .RESET_B(_00516_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[72] ));
 sky130_fd_sc_hd__dfrtp_2 _11127_ (.CLK(clknet_leaf_62_clk),
    .D(_01692_),
    .RESET_B(_00517_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[73] ));
 sky130_fd_sc_hd__dfrtp_2 _11128_ (.CLK(clknet_leaf_59_clk),
    .D(_01693_),
    .RESET_B(_00518_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[74] ));
 sky130_fd_sc_hd__dfrtp_2 _11129_ (.CLK(clknet_leaf_60_clk),
    .D(_01694_),
    .RESET_B(_00519_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[75] ));
 sky130_fd_sc_hd__dfrtp_2 _11130_ (.CLK(clknet_leaf_59_clk),
    .D(_01695_),
    .RESET_B(_00520_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[76] ));
 sky130_fd_sc_hd__dfrtp_1 _11131_ (.CLK(clknet_leaf_60_clk),
    .D(_01696_),
    .RESET_B(_00521_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[77] ));
 sky130_fd_sc_hd__dfrtp_1 _11132_ (.CLK(clknet_leaf_59_clk),
    .D(_01697_),
    .RESET_B(_00522_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[78] ));
 sky130_fd_sc_hd__dfrtp_1 _11133_ (.CLK(clknet_leaf_58_clk),
    .D(_01698_),
    .RESET_B(_00523_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[79] ));
 sky130_fd_sc_hd__dfrtp_2 _11134_ (.CLK(clknet_leaf_58_clk),
    .D(_01699_),
    .RESET_B(_00524_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[80] ));
 sky130_fd_sc_hd__dfrtp_2 _11135_ (.CLK(clknet_leaf_58_clk),
    .D(_01700_),
    .RESET_B(_00525_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[81] ));
 sky130_fd_sc_hd__dfrtp_2 _11136_ (.CLK(clknet_leaf_54_clk),
    .D(_01701_),
    .RESET_B(_00526_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[82] ));
 sky130_fd_sc_hd__dfrtp_2 _11137_ (.CLK(clknet_leaf_54_clk),
    .D(_01702_),
    .RESET_B(_00527_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[83] ));
 sky130_fd_sc_hd__dfrtp_2 _11138_ (.CLK(clknet_leaf_54_clk),
    .D(_01703_),
    .RESET_B(_00528_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[84] ));
 sky130_fd_sc_hd__dfrtp_1 _11139_ (.CLK(clknet_leaf_53_clk),
    .D(_01704_),
    .RESET_B(_00529_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[85] ));
 sky130_fd_sc_hd__dfrtp_1 _11140_ (.CLK(clknet_leaf_53_clk),
    .D(_01705_),
    .RESET_B(_00530_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[86] ));
 sky130_fd_sc_hd__dfrtp_2 _11141_ (.CLK(clknet_leaf_53_clk),
    .D(_01706_),
    .RESET_B(_00531_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[87] ));
 sky130_fd_sc_hd__dfrtp_2 _11142_ (.CLK(clknet_leaf_52_clk),
    .D(_01707_),
    .RESET_B(_00532_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[88] ));
 sky130_fd_sc_hd__dfrtp_2 _11143_ (.CLK(clknet_leaf_36_clk),
    .D(_01708_),
    .RESET_B(_00533_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[89] ));
 sky130_fd_sc_hd__dfrtp_1 _11144_ (.CLK(clknet_leaf_35_clk),
    .D(_01709_),
    .RESET_B(_00534_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[90] ));
 sky130_fd_sc_hd__dfrtp_2 _11145_ (.CLK(clknet_leaf_35_clk),
    .D(_01710_),
    .RESET_B(_00535_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[91] ));
 sky130_fd_sc_hd__dfrtp_2 _11146_ (.CLK(clknet_leaf_34_clk),
    .D(_01711_),
    .RESET_B(_00536_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[92] ));
 sky130_fd_sc_hd__dfrtp_2 _11147_ (.CLK(clknet_leaf_34_clk),
    .D(_01712_),
    .RESET_B(_00537_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[93] ));
 sky130_fd_sc_hd__dfrtp_2 _11148_ (.CLK(clknet_leaf_35_clk),
    .D(_01713_),
    .RESET_B(_00538_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[94] ));
 sky130_fd_sc_hd__dfrtp_2 _11149_ (.CLK(clknet_leaf_35_clk),
    .D(_01714_),
    .RESET_B(_00539_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[95] ));
 sky130_fd_sc_hd__dfrtp_4 _11150_ (.CLK(clknet_leaf_40_clk),
    .D(_01715_),
    .RESET_B(_00540_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[96] ));
 sky130_fd_sc_hd__dfrtp_4 _11151_ (.CLK(clknet_leaf_46_clk),
    .D(_01716_),
    .RESET_B(_00541_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[97] ));
 sky130_fd_sc_hd__dfrtp_4 _11152_ (.CLK(clknet_leaf_64_clk),
    .D(_01717_),
    .RESET_B(_00542_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[98] ));
 sky130_fd_sc_hd__dfrtp_1 _11153_ (.CLK(clknet_leaf_63_clk),
    .D(_01718_),
    .RESET_B(_00543_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[99] ));
 sky130_fd_sc_hd__dfrtp_2 _11154_ (.CLK(clknet_leaf_63_clk),
    .D(_01719_),
    .RESET_B(_00544_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[100] ));
 sky130_fd_sc_hd__dfrtp_1 _11155_ (.CLK(clknet_leaf_64_clk),
    .D(_01720_),
    .RESET_B(_00545_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[101] ));
 sky130_fd_sc_hd__dfrtp_1 _11156_ (.CLK(clknet_leaf_64_clk),
    .D(_01721_),
    .RESET_B(_00546_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[102] ));
 sky130_fd_sc_hd__dfrtp_2 _11157_ (.CLK(clknet_leaf_64_clk),
    .D(_01722_),
    .RESET_B(_00547_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[103] ));
 sky130_fd_sc_hd__dfrtp_2 _11158_ (.CLK(clknet_leaf_64_clk),
    .D(_01723_),
    .RESET_B(_00548_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[104] ));
 sky130_fd_sc_hd__dfrtp_2 _11159_ (.CLK(clknet_leaf_62_clk),
    .D(_01724_),
    .RESET_B(_00549_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[105] ));
 sky130_fd_sc_hd__dfrtp_2 _11160_ (.CLK(clknet_leaf_60_clk),
    .D(_01725_),
    .RESET_B(_00550_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[106] ));
 sky130_fd_sc_hd__dfrtp_2 _11161_ (.CLK(clknet_leaf_61_clk),
    .D(_01726_),
    .RESET_B(_00551_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[107] ));
 sky130_fd_sc_hd__dfrtp_2 _11162_ (.CLK(clknet_leaf_60_clk),
    .D(_01727_),
    .RESET_B(_00552_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[108] ));
 sky130_fd_sc_hd__dfrtp_1 _11163_ (.CLK(clknet_leaf_60_clk),
    .D(_01728_),
    .RESET_B(_00553_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[109] ));
 sky130_fd_sc_hd__dfrtp_1 _11164_ (.CLK(clknet_leaf_59_clk),
    .D(_01729_),
    .RESET_B(_00554_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[110] ));
 sky130_fd_sc_hd__dfrtp_2 _11165_ (.CLK(clknet_leaf_57_clk),
    .D(_01730_),
    .RESET_B(_00555_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[111] ));
 sky130_fd_sc_hd__dfrtp_2 _11166_ (.CLK(clknet_leaf_57_clk),
    .D(_01731_),
    .RESET_B(_00556_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[112] ));
 sky130_fd_sc_hd__dfrtp_2 _11167_ (.CLK(clknet_leaf_54_clk),
    .D(_01732_),
    .RESET_B(_00557_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[113] ));
 sky130_fd_sc_hd__dfrtp_2 _11168_ (.CLK(clknet_leaf_54_clk),
    .D(_01733_),
    .RESET_B(_00558_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[114] ));
 sky130_fd_sc_hd__dfrtp_1 _11169_ (.CLK(clknet_leaf_55_clk),
    .D(_01734_),
    .RESET_B(_00559_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[115] ));
 sky130_fd_sc_hd__dfrtp_1 _11170_ (.CLK(clknet_leaf_55_clk),
    .D(_01735_),
    .RESET_B(_00560_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[116] ));
 sky130_fd_sc_hd__dfrtp_2 _11171_ (.CLK(clknet_leaf_49_clk),
    .D(_01736_),
    .RESET_B(_00561_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[117] ));
 sky130_fd_sc_hd__dfrtp_1 _11172_ (.CLK(clknet_leaf_49_clk),
    .D(_01737_),
    .RESET_B(_00562_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[118] ));
 sky130_fd_sc_hd__dfrtp_2 _11173_ (.CLK(clknet_leaf_51_clk),
    .D(_01738_),
    .RESET_B(_00563_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[119] ));
 sky130_fd_sc_hd__dfrtp_2 _11174_ (.CLK(clknet_leaf_37_clk),
    .D(_01739_),
    .RESET_B(_00564_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[120] ));
 sky130_fd_sc_hd__dfrtp_1 _11175_ (.CLK(clknet_leaf_37_clk),
    .D(_01740_),
    .RESET_B(_00565_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[121] ));
 sky130_fd_sc_hd__dfrtp_1 _11176_ (.CLK(clknet_leaf_37_clk),
    .D(_01741_),
    .RESET_B(_00566_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[122] ));
 sky130_fd_sc_hd__dfrtp_1 _11177_ (.CLK(clknet_leaf_35_clk),
    .D(_01742_),
    .RESET_B(_00567_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[123] ));
 sky130_fd_sc_hd__dfrtp_2 _11178_ (.CLK(clknet_leaf_38_clk),
    .D(_01743_),
    .RESET_B(_00568_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[124] ));
 sky130_fd_sc_hd__dfrtp_1 _11179_ (.CLK(clknet_leaf_38_clk),
    .D(_01744_),
    .RESET_B(_00569_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[125] ));
 sky130_fd_sc_hd__dfrtp_2 _11180_ (.CLK(clknet_leaf_38_clk),
    .D(_01745_),
    .RESET_B(_00570_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[126] ));
 sky130_fd_sc_hd__dfrtp_1 _11181_ (.CLK(clknet_leaf_33_clk),
    .D(_01746_),
    .RESET_B(_00571_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.char_path_n[127] ));
 sky130_fd_sc_hd__dfrtp_1 _11182_ (.CLK(clknet_leaf_33_clk),
    .D(_01747_),
    .RESET_B(_00572_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.curr_path[127] ));
 sky130_fd_sc_hd__dfrtp_4 _11183_ (.CLK(clknet_leaf_34_clk),
    .D(_01748_),
    .RESET_B(_00573_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.cb_length[0] ));
 sky130_fd_sc_hd__dfrtp_2 _11184_ (.CLK(clknet_leaf_34_clk),
    .D(_01749_),
    .RESET_B(_00574_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.cb_length[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11185_ (.CLK(clknet_leaf_34_clk),
    .D(_01750_),
    .RESET_B(_00575_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.cb_length[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11186_ (.CLK(clknet_leaf_34_clk),
    .D(_01751_),
    .RESET_B(_00576_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.cb_length[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11187_ (.CLK(clknet_leaf_33_clk),
    .D(_01752_),
    .RESET_B(_00577_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.cb_length[4] ));
 sky130_fd_sc_hd__dfrtp_1 _11188_ (.CLK(clknet_leaf_33_clk),
    .D(_01753_),
    .RESET_B(_00578_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.cb_length[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11189_ (.CLK(clknet_leaf_33_clk),
    .D(_01754_),
    .RESET_B(_00579_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.cb_length[6] ));
 sky130_fd_sc_hd__dfrtp_1 _11190_ (.CLK(clknet_leaf_27_clk),
    .D(_01755_),
    .RESET_B(_00580_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.num_lefts[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11191_ (.CLK(clknet_leaf_27_clk),
    .D(_01756_),
    .RESET_B(_00581_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.num_lefts[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11192_ (.CLK(clknet_leaf_27_clk),
    .D(_01757_),
    .RESET_B(_00582_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.num_lefts[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11193_ (.CLK(clknet_leaf_27_clk),
    .D(_01758_),
    .RESET_B(_00583_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.num_lefts[3] ));
 sky130_fd_sc_hd__dfrtp_2 _11194_ (.CLK(clknet_leaf_27_clk),
    .D(_01759_),
    .RESET_B(_00584_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.num_lefts[4] ));
 sky130_fd_sc_hd__dfrtp_1 _11195_ (.CLK(clknet_leaf_28_clk),
    .D(_01760_),
    .RESET_B(_00585_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.num_lefts[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11196_ (.CLK(clknet_leaf_26_clk),
    .D(_01761_),
    .RESET_B(_00586_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.num_lefts[6] ));
 sky130_fd_sc_hd__dfrtp_1 _11197_ (.CLK(clknet_leaf_26_clk),
    .D(_01762_),
    .RESET_B(_00587_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.num_lefts[7] ));
 sky130_fd_sc_hd__dfrtp_1 _11198_ (.CLK(clknet_leaf_32_clk),
    .D(_01763_),
    .RESET_B(_00588_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.left ));
 sky130_fd_sc_hd__dfrtp_2 _11199_ (.CLK(clknet_leaf_29_clk),
    .D(_01764_),
    .RESET_B(_00589_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.zeroes[0] ));
 sky130_fd_sc_hd__dfrtp_2 _11200_ (.CLK(clknet_leaf_30_clk),
    .D(_01765_),
    .RESET_B(_00590_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.zeroes[1] ));
 sky130_fd_sc_hd__dfrtp_2 _11201_ (.CLK(clknet_leaf_29_clk),
    .D(_01766_),
    .RESET_B(_00591_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.zeroes[2] ));
 sky130_fd_sc_hd__dfrtp_2 _11202_ (.CLK(clknet_leaf_30_clk),
    .D(_01767_),
    .RESET_B(_00592_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.zeroes[3] ));
 sky130_fd_sc_hd__dfrtp_2 _11203_ (.CLK(clknet_leaf_30_clk),
    .D(_01768_),
    .RESET_B(_00593_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.zeroes[4] ));
 sky130_fd_sc_hd__dfrtp_1 _11204_ (.CLK(clknet_leaf_30_clk),
    .D(_01769_),
    .RESET_B(_00594_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.zeroes[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11205_ (.CLK(clknet_leaf_30_clk),
    .D(_01770_),
    .RESET_B(_00595_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.zeroes[6] ));
 sky130_fd_sc_hd__dfrtp_1 _11206_ (.CLK(clknet_leaf_26_clk),
    .D(_01771_),
    .RESET_B(_00596_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.zeroes[7] ));
 sky130_fd_sc_hd__dfstp_1 _11207_ (.CLK(clknet_leaf_26_clk),
    .D(_01772_),
    .SET_B(_00597_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.wait_cycle ));
 sky130_fd_sc_hd__dfstp_1 _11208_ (.CLK(clknet_leaf_25_clk),
    .D(_01773_),
    .SET_B(_00598_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.setup ));
 sky130_fd_sc_hd__dfrtp_2 _11209_ (.CLK(clknet_leaf_107_clk),
    .D(_01774_),
    .RESET_B(_00599_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.alternator_timer[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11210_ (.CLK(clknet_leaf_107_clk),
    .D(_01775_),
    .RESET_B(_00600_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.alternator_timer[1] ));
 sky130_fd_sc_hd__dfrtp_2 _11211_ (.CLK(clknet_leaf_107_clk),
    .D(_01776_),
    .RESET_B(_00601_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.alternator_timer[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11212_ (.CLK(clknet_leaf_107_clk),
    .D(_01777_),
    .RESET_B(_00602_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.alternator_timer[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11213_ (.CLK(clknet_leaf_105_clk),
    .D(_01778_),
    .RESET_B(_00603_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.wait_cnt ));
 sky130_fd_sc_hd__dfrtp_1 _11214_ (.CLK(clknet_leaf_15_clk),
    .D(_01779_),
    .RESET_B(_00604_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.nullSumIndex[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11215_ (.CLK(clknet_leaf_43_clk),
    .D(_01780_),
    .RESET_B(_00605_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.nullSumIndex[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11216_ (.CLK(clknet_leaf_15_clk),
    .D(_01781_),
    .RESET_B(_00606_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.nullSumIndex[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11217_ (.CLK(clknet_leaf_14_clk),
    .D(_01782_),
    .RESET_B(_00607_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.nullSumIndex[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11218_ (.CLK(clknet_leaf_14_clk),
    .D(_01783_),
    .RESET_B(_00608_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.nullSumIndex[4] ));
 sky130_fd_sc_hd__dfrtp_1 _11219_ (.CLK(clknet_leaf_43_clk),
    .D(_01784_),
    .RESET_B(_00609_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.nullSumIndex[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11220_ (.CLK(clknet_leaf_43_clk),
    .D(_01785_),
    .RESET_B(_00610_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.nullSumIndex[6] ));
 sky130_fd_sc_hd__dfrtp_1 _11221_ (.CLK(clknet_leaf_106_clk),
    .D(net1005),
    .RESET_B(_00611_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.HT_fin_reg ));
 sky130_fd_sc_hd__dfrtp_1 _11222_ (.CLK(clknet_leaf_106_clk),
    .D(_01787_),
    .RESET_B(_00612_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.controller.fin_FINISHED ));
 sky130_fd_sc_hd__dfrtp_4 _11223_ (.CLK(clknet_leaf_12_clk),
    .D(_01788_),
    .RESET_B(_00613_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.WorR ));
 sky130_fd_sc_hd__dfrtp_1 _11224_ (.CLK(clknet_leaf_83_clk),
    .D(_01789_),
    .RESET_B(_00614_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11225_ (.CLK(clknet_leaf_85_clk),
    .D(_01790_),
    .RESET_B(_00615_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11226_ (.CLK(clknet_leaf_83_clk),
    .D(_01791_),
    .RESET_B(_00616_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11227_ (.CLK(clknet_leaf_84_clk),
    .D(_01792_),
    .RESET_B(_00617_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11228_ (.CLK(clknet_leaf_84_clk),
    .D(_01793_),
    .RESET_B(_00618_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[4] ));
 sky130_fd_sc_hd__dfrtp_1 _11229_ (.CLK(clknet_leaf_83_clk),
    .D(_01794_),
    .RESET_B(_00619_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11230_ (.CLK(clknet_leaf_82_clk),
    .D(_01795_),
    .RESET_B(_00620_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[6] ));
 sky130_fd_sc_hd__dfrtp_1 _11231_ (.CLK(clknet_leaf_83_clk),
    .D(_01796_),
    .RESET_B(_00621_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[7] ));
 sky130_fd_sc_hd__dfrtp_1 _11232_ (.CLK(clknet_leaf_66_clk),
    .D(_01797_),
    .RESET_B(_00622_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[8] ));
 sky130_fd_sc_hd__dfrtp_1 _11233_ (.CLK(clknet_leaf_82_clk),
    .D(_01798_),
    .RESET_B(_00623_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[9] ));
 sky130_fd_sc_hd__dfrtp_1 _11234_ (.CLK(clknet_leaf_82_clk),
    .D(net1590),
    .RESET_B(_00624_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[10] ));
 sky130_fd_sc_hd__dfrtp_1 _11235_ (.CLK(clknet_leaf_67_clk),
    .D(net1601),
    .RESET_B(_00625_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[11] ));
 sky130_fd_sc_hd__dfrtp_1 _11236_ (.CLK(clknet_leaf_66_clk),
    .D(_01801_),
    .RESET_B(_00626_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[12] ));
 sky130_fd_sc_hd__dfrtp_1 _11237_ (.CLK(clknet_leaf_67_clk),
    .D(net1560),
    .RESET_B(_00627_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[13] ));
 sky130_fd_sc_hd__dfrtp_1 _11238_ (.CLK(clknet_leaf_67_clk),
    .D(_01803_),
    .RESET_B(_00628_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[14] ));
 sky130_fd_sc_hd__dfrtp_1 _11239_ (.CLK(clknet_leaf_67_clk),
    .D(net1437),
    .RESET_B(_00629_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[15] ));
 sky130_fd_sc_hd__dfrtp_1 _11240_ (.CLK(clknet_leaf_69_clk),
    .D(net1568),
    .RESET_B(_00630_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[16] ));
 sky130_fd_sc_hd__dfrtp_1 _11241_ (.CLK(clknet_leaf_69_clk),
    .D(net1444),
    .RESET_B(_00631_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[17] ));
 sky130_fd_sc_hd__dfrtp_1 _11242_ (.CLK(clknet_leaf_69_clk),
    .D(net1571),
    .RESET_B(_00632_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[18] ));
 sky130_fd_sc_hd__dfrtp_1 _11243_ (.CLK(clknet_leaf_77_clk),
    .D(net1351),
    .RESET_B(_00633_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[19] ));
 sky130_fd_sc_hd__dfrtp_1 _11244_ (.CLK(clknet_leaf_77_clk),
    .D(net1396),
    .RESET_B(_00634_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[20] ));
 sky130_fd_sc_hd__dfrtp_1 _11245_ (.CLK(clknet_leaf_73_clk),
    .D(net1553),
    .RESET_B(_00635_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[21] ));
 sky130_fd_sc_hd__dfrtp_1 _11246_ (.CLK(clknet_leaf_73_clk),
    .D(_01811_),
    .RESET_B(_00636_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[22] ));
 sky130_fd_sc_hd__dfrtp_1 _11247_ (.CLK(clknet_leaf_77_clk),
    .D(_01812_),
    .RESET_B(_00637_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[23] ));
 sky130_fd_sc_hd__dfrtp_1 _11248_ (.CLK(clknet_leaf_76_clk),
    .D(net1432),
    .RESET_B(_00638_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[24] ));
 sky130_fd_sc_hd__dfrtp_1 _11249_ (.CLK(clknet_leaf_74_clk),
    .D(net1566),
    .RESET_B(_00639_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[25] ));
 sky130_fd_sc_hd__dfrtp_1 _11250_ (.CLK(clknet_leaf_75_clk),
    .D(net1547),
    .RESET_B(_00640_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[26] ));
 sky130_fd_sc_hd__dfrtp_1 _11251_ (.CLK(clknet_leaf_76_clk),
    .D(_01816_),
    .RESET_B(_00641_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[27] ));
 sky130_fd_sc_hd__dfrtp_1 _11252_ (.CLK(clknet_leaf_103_clk),
    .D(_01817_),
    .RESET_B(_00642_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[28] ));
 sky130_fd_sc_hd__dfrtp_1 _11253_ (.CLK(clknet_leaf_106_clk),
    .D(net1494),
    .RESET_B(_00643_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[29] ));
 sky130_fd_sc_hd__dfrtp_1 _11254_ (.CLK(clknet_leaf_103_clk),
    .D(net1491),
    .RESET_B(_00644_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[30] ));
 sky130_fd_sc_hd__dfrtp_1 _11255_ (.CLK(clknet_leaf_105_clk),
    .D(_01820_),
    .RESET_B(_00645_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[31] ));
 sky130_fd_sc_hd__dfrtp_1 _11256_ (.CLK(clknet_leaf_79_clk),
    .D(_01821_),
    .RESET_B(_00646_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[32] ));
 sky130_fd_sc_hd__dfrtp_1 _11257_ (.CLK(clknet_leaf_80_clk),
    .D(net1586),
    .RESET_B(_00647_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[33] ));
 sky130_fd_sc_hd__dfrtp_1 _11258_ (.CLK(clknet_leaf_79_clk),
    .D(_01823_),
    .RESET_B(_00648_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[34] ));
 sky130_fd_sc_hd__dfrtp_1 _11259_ (.CLK(clknet_leaf_80_clk),
    .D(_01824_),
    .RESET_B(_00649_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[35] ));
 sky130_fd_sc_hd__dfrtp_1 _11260_ (.CLK(clknet_leaf_80_clk),
    .D(_01825_),
    .RESET_B(_00650_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[36] ));
 sky130_fd_sc_hd__dfrtp_1 _11261_ (.CLK(clknet_leaf_81_clk),
    .D(_01826_),
    .RESET_B(_00651_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[37] ));
 sky130_fd_sc_hd__dfrtp_1 _11262_ (.CLK(clknet_leaf_81_clk),
    .D(_01827_),
    .RESET_B(_00652_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[38] ));
 sky130_fd_sc_hd__dfrtp_1 _11263_ (.CLK(clknet_leaf_81_clk),
    .D(_01828_),
    .RESET_B(_00653_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[39] ));
 sky130_fd_sc_hd__dfrtp_1 _11264_ (.CLK(clknet_leaf_68_clk),
    .D(_01829_),
    .RESET_B(_00654_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[40] ));
 sky130_fd_sc_hd__dfrtp_1 _11265_ (.CLK(clknet_leaf_81_clk),
    .D(_01830_),
    .RESET_B(_00655_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[41] ));
 sky130_fd_sc_hd__dfrtp_1 _11266_ (.CLK(clknet_leaf_82_clk),
    .D(_01831_),
    .RESET_B(_00656_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[42] ));
 sky130_fd_sc_hd__dfrtp_1 _11267_ (.CLK(clknet_leaf_68_clk),
    .D(_01832_),
    .RESET_B(_00657_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[43] ));
 sky130_fd_sc_hd__dfrtp_1 _11268_ (.CLK(clknet_leaf_69_clk),
    .D(net1451),
    .RESET_B(_00658_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[44] ));
 sky130_fd_sc_hd__dfrtp_1 _11269_ (.CLK(clknet_leaf_69_clk),
    .D(_01834_),
    .RESET_B(_00659_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[45] ));
 sky130_fd_sc_hd__dfrtp_1 _11270_ (.CLK(clknet_leaf_45_clk),
    .D(_01835_),
    .RESET_B(_00660_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[46] ));
 sky130_fd_sc_hd__dfrtp_1 _11271_ (.CLK(clknet_leaf_43_clk),
    .D(_01836_),
    .RESET_B(_00661_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[47] ));
 sky130_fd_sc_hd__dfrtp_1 _11272_ (.CLK(clknet_leaf_42_clk),
    .D(_01837_),
    .RESET_B(_00662_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[48] ));
 sky130_fd_sc_hd__dfrtp_1 _11273_ (.CLK(clknet_leaf_44_clk),
    .D(_01838_),
    .RESET_B(_00663_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[49] ));
 sky130_fd_sc_hd__dfrtp_1 _11274_ (.CLK(clknet_leaf_44_clk),
    .D(_01839_),
    .RESET_B(_00664_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[50] ));
 sky130_fd_sc_hd__dfrtp_1 _11275_ (.CLK(clknet_leaf_42_clk),
    .D(_01840_),
    .RESET_B(_00665_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[51] ));
 sky130_fd_sc_hd__dfrtp_1 _11276_ (.CLK(clknet_leaf_43_clk),
    .D(_01841_),
    .RESET_B(_00666_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[52] ));
 sky130_fd_sc_hd__dfrtp_1 _11277_ (.CLK(clknet_leaf_44_clk),
    .D(_01842_),
    .RESET_B(_00667_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[53] ));
 sky130_fd_sc_hd__dfrtp_1 _11278_ (.CLK(clknet_leaf_104_clk),
    .D(_01843_),
    .RESET_B(_00668_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[54] ));
 sky130_fd_sc_hd__dfrtp_1 _11279_ (.CLK(clknet_leaf_44_clk),
    .D(_01844_),
    .RESET_B(_00669_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[55] ));
 sky130_fd_sc_hd__dfrtp_1 _11280_ (.CLK(clknet_leaf_45_clk),
    .D(_01845_),
    .RESET_B(_00670_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[56] ));
 sky130_fd_sc_hd__dfrtp_1 _11281_ (.CLK(clknet_leaf_44_clk),
    .D(_01846_),
    .RESET_B(_00671_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[57] ));
 sky130_fd_sc_hd__dfrtp_1 _11282_ (.CLK(clknet_leaf_44_clk),
    .D(_01847_),
    .RESET_B(_00672_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[58] ));
 sky130_fd_sc_hd__dfrtp_1 _11283_ (.CLK(clknet_leaf_44_clk),
    .D(_01848_),
    .RESET_B(_00673_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[59] ));
 sky130_fd_sc_hd__dfrtp_1 _11284_ (.CLK(clknet_leaf_42_clk),
    .D(_01849_),
    .RESET_B(_00674_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[60] ));
 sky130_fd_sc_hd__dfrtp_1 _11285_ (.CLK(clknet_leaf_44_clk),
    .D(_01850_),
    .RESET_B(_00675_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[61] ));
 sky130_fd_sc_hd__dfrtp_1 _11286_ (.CLK(clknet_leaf_14_clk),
    .D(_01851_),
    .RESET_B(_00676_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[62] ));
 sky130_fd_sc_hd__dfrtp_1 _11287_ (.CLK(clknet_leaf_104_clk),
    .D(_01852_),
    .RESET_B(_00677_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.tree_reg[63] ));
 sky130_fd_sc_hd__dfrtp_1 _11288_ (.CLK(clknet_leaf_14_clk),
    .D(_01853_),
    .RESET_B(_00678_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.closing ));
 sky130_fd_sc_hd__dfrtp_1 _11289_ (.CLK(clknet_leaf_24_clk),
    .D(_01854_),
    .RESET_B(_00679_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.curr_index[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11290_ (.CLK(clknet_leaf_20_clk),
    .D(_01855_),
    .RESET_B(_00680_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.curr_index[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11291_ (.CLK(clknet_leaf_22_clk),
    .D(_01856_),
    .RESET_B(_00681_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.curr_index[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11292_ (.CLK(clknet_leaf_24_clk),
    .D(_01857_),
    .RESET_B(_00682_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.curr_index[4] ));
 sky130_fd_sc_hd__dfrtp_1 _11293_ (.CLK(clknet_leaf_24_clk),
    .D(_01858_),
    .RESET_B(_00683_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.curr_index[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11294_ (.CLK(clknet_leaf_22_clk),
    .D(_01859_),
    .RESET_B(_00684_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.curr_index[6] ));
 sky130_fd_sc_hd__dfrtp_1 _11295_ (.CLK(clknet_leaf_24_clk),
    .D(_01860_),
    .RESET_B(_00685_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.curr_index[7] ));
 sky130_fd_sc_hd__dfrtp_1 _11296_ (.CLK(clknet_leaf_2_clk),
    .D(_01861_),
    .RESET_B(_00686_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.dut.out[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11297_ (.CLK(clknet_leaf_2_clk),
    .D(_01862_),
    .RESET_B(_00687_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.dut.out[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11298_ (.CLK(clknet_leaf_5_clk),
    .D(_01863_),
    .RESET_B(_00688_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.dut.out[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11299_ (.CLK(clknet_leaf_4_clk),
    .D(_01864_),
    .RESET_B(_00689_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.dut.out[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11300_ (.CLK(clknet_leaf_2_clk),
    .D(_01865_),
    .RESET_B(_00690_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.dut.out[4] ));
 sky130_fd_sc_hd__dfrtp_1 _11301_ (.CLK(clknet_leaf_2_clk),
    .D(_01866_),
    .RESET_B(_00691_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.dut.out[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11302_ (.CLK(clknet_leaf_2_clk),
    .D(_01867_),
    .RESET_B(_00692_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.dut.out[6] ));
 sky130_fd_sc_hd__dfrtp_1 _11303_ (.CLK(clknet_leaf_0_clk),
    .D(_01868_),
    .RESET_B(_00693_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.dut.out[7] ));
 sky130_fd_sc_hd__dfrtp_2 _11304_ (.CLK(clknet_leaf_43_clk),
    .D(_01869_),
    .RESET_B(_00694_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.least1[0] ));
 sky130_fd_sc_hd__dfrtp_2 _11305_ (.CLK(clknet_leaf_43_clk),
    .D(_01870_),
    .RESET_B(_00695_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.least1[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11306_ (.CLK(clknet_leaf_43_clk),
    .D(_01871_),
    .RESET_B(_00696_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.least1[2] ));
 sky130_fd_sc_hd__dfrtp_2 _11307_ (.CLK(clknet_leaf_43_clk),
    .D(_01872_),
    .RESET_B(_00697_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.least1[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11308_ (.CLK(clknet_leaf_14_clk),
    .D(_01873_),
    .RESET_B(_00698_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.least1[4] ));
 sky130_fd_sc_hd__dfrtp_2 _11309_ (.CLK(clknet_leaf_14_clk),
    .D(_01874_),
    .RESET_B(_00699_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.least1[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11310_ (.CLK(clknet_leaf_43_clk),
    .D(_01875_),
    .RESET_B(_00700_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.least1[6] ));
 sky130_fd_sc_hd__dfstp_1 _11311_ (.CLK(clknet_leaf_14_clk),
    .D(_01876_),
    .SET_B(_00701_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.least1[7] ));
 sky130_fd_sc_hd__dfstp_1 _11312_ (.CLK(clknet_leaf_13_clk),
    .D(_01877_),
    .SET_B(_00702_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.least1[8] ));
 sky130_fd_sc_hd__dfrtp_2 _11313_ (.CLK(clknet_leaf_41_clk),
    .D(_01878_),
    .RESET_B(_00703_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.least2[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11314_ (.CLK(clknet_leaf_41_clk),
    .D(_01879_),
    .RESET_B(_00704_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.least2[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11315_ (.CLK(clknet_leaf_43_clk),
    .D(_01880_),
    .RESET_B(_00705_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.least2[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11316_ (.CLK(clknet_leaf_44_clk),
    .D(_01881_),
    .RESET_B(_00706_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.least2[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11317_ (.CLK(clknet_leaf_44_clk),
    .D(_01882_),
    .RESET_B(_00707_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.least2[4] ));
 sky130_fd_sc_hd__dfrtp_1 _11318_ (.CLK(clknet_leaf_41_clk),
    .D(_01883_),
    .RESET_B(_00708_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.least2[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11319_ (.CLK(clknet_leaf_43_clk),
    .D(_01884_),
    .RESET_B(_00709_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.least2[6] ));
 sky130_fd_sc_hd__dfstp_1 _11320_ (.CLK(clknet_leaf_14_clk),
    .D(_01885_),
    .SET_B(_00710_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.least2[7] ));
 sky130_fd_sc_hd__dfstp_2 _11321_ (.CLK(clknet_leaf_104_clk),
    .D(_01886_),
    .SET_B(_00711_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.least2[8] ));
 sky130_fd_sc_hd__dfrtp_2 _11322_ (.CLK(clknet_leaf_90_clk),
    .D(_01887_),
    .RESET_B(_00712_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.sum[0] ));
 sky130_fd_sc_hd__dfrtp_2 _11323_ (.CLK(clknet_leaf_90_clk),
    .D(_01888_),
    .RESET_B(_00713_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.sum[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11324_ (.CLK(clknet_leaf_89_clk),
    .D(_01889_),
    .RESET_B(_00714_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.sum[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11325_ (.CLK(clknet_leaf_89_clk),
    .D(_01890_),
    .RESET_B(_00715_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.sum[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11326_ (.CLK(clknet_leaf_88_clk),
    .D(_01891_),
    .RESET_B(_00716_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.sum[4] ));
 sky130_fd_sc_hd__dfrtp_1 _11327_ (.CLK(clknet_leaf_88_clk),
    .D(_01892_),
    .RESET_B(_00717_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.sum[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11328_ (.CLK(clknet_leaf_88_clk),
    .D(_01893_),
    .RESET_B(_00718_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.sum[6] ));
 sky130_fd_sc_hd__dfrtp_1 _11329_ (.CLK(clknet_leaf_88_clk),
    .D(_01894_),
    .RESET_B(_00719_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.sum[7] ));
 sky130_fd_sc_hd__dfrtp_1 _11330_ (.CLK(clknet_leaf_82_clk),
    .D(_01895_),
    .RESET_B(_00720_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.sum[8] ));
 sky130_fd_sc_hd__dfrtp_1 _11331_ (.CLK(clknet_leaf_84_clk),
    .D(_01896_),
    .RESET_B(_00721_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.sum[9] ));
 sky130_fd_sc_hd__dfrtp_1 _11332_ (.CLK(clknet_leaf_84_clk),
    .D(_01897_),
    .RESET_B(_00722_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.sum[10] ));
 sky130_fd_sc_hd__dfrtp_1 _11333_ (.CLK(clknet_leaf_84_clk),
    .D(_01898_),
    .RESET_B(_00723_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.sum[11] ));
 sky130_fd_sc_hd__dfrtp_1 _11334_ (.CLK(clknet_leaf_82_clk),
    .D(_01899_),
    .RESET_B(_00724_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.sum[12] ));
 sky130_fd_sc_hd__dfrtp_2 _11335_ (.CLK(clknet_leaf_84_clk),
    .D(_01900_),
    .RESET_B(_00725_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.sum[13] ));
 sky130_fd_sc_hd__dfrtp_1 _11336_ (.CLK(clknet_leaf_81_clk),
    .D(_01901_),
    .RESET_B(_00726_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.sum[14] ));
 sky130_fd_sc_hd__dfrtp_1 _11337_ (.CLK(clknet_leaf_84_clk),
    .D(_01902_),
    .RESET_B(_00727_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.sum[15] ));
 sky130_fd_sc_hd__dfrtp_1 _11338_ (.CLK(clknet_leaf_77_clk),
    .D(_01903_),
    .RESET_B(_00728_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.sum[16] ));
 sky130_fd_sc_hd__dfrtp_1 _11339_ (.CLK(clknet_leaf_77_clk),
    .D(_01904_),
    .RESET_B(_00729_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.sum[17] ));
 sky130_fd_sc_hd__dfrtp_1 _11340_ (.CLK(clknet_leaf_77_clk),
    .D(_01905_),
    .RESET_B(_00730_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.sum[18] ));
 sky130_fd_sc_hd__dfrtp_1 _11341_ (.CLK(clknet_leaf_77_clk),
    .D(_01906_),
    .RESET_B(_00731_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.sum[19] ));
 sky130_fd_sc_hd__dfrtp_1 _11342_ (.CLK(clknet_leaf_77_clk),
    .D(_01907_),
    .RESET_B(_00732_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.sum[20] ));
 sky130_fd_sc_hd__dfrtp_1 _11343_ (.CLK(clknet_leaf_77_clk),
    .D(_01908_),
    .RESET_B(_00733_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.sum[21] ));
 sky130_fd_sc_hd__dfrtp_1 _11344_ (.CLK(clknet_leaf_76_clk),
    .D(_01909_),
    .RESET_B(_00734_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.sum[22] ));
 sky130_fd_sc_hd__dfrtp_1 _11345_ (.CLK(clknet_leaf_76_clk),
    .D(_01910_),
    .RESET_B(_00735_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.sum[23] ));
 sky130_fd_sc_hd__dfrtp_1 _11346_ (.CLK(clknet_leaf_76_clk),
    .D(_01911_),
    .RESET_B(_00736_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.sum[24] ));
 sky130_fd_sc_hd__dfrtp_1 _11347_ (.CLK(clknet_leaf_76_clk),
    .D(_01912_),
    .RESET_B(_00737_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.sum[25] ));
 sky130_fd_sc_hd__dfrtp_1 _11348_ (.CLK(clknet_leaf_75_clk),
    .D(_01913_),
    .RESET_B(_00738_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.sum[26] ));
 sky130_fd_sc_hd__dfrtp_1 _11349_ (.CLK(clknet_leaf_103_clk),
    .D(_01914_),
    .RESET_B(_00739_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.sum[27] ));
 sky130_fd_sc_hd__dfrtp_1 _11350_ (.CLK(clknet_leaf_103_clk),
    .D(_01915_),
    .RESET_B(_00740_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.sum[28] ));
 sky130_fd_sc_hd__dfrtp_1 _11351_ (.CLK(clknet_leaf_106_clk),
    .D(_01916_),
    .RESET_B(_00741_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.sum[29] ));
 sky130_fd_sc_hd__dfrtp_1 _11352_ (.CLK(clknet_leaf_103_clk),
    .D(_01917_),
    .RESET_B(_00742_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.sum[30] ));
 sky130_fd_sc_hd__dfrtp_1 _11353_ (.CLK(clknet_leaf_106_clk),
    .D(_01918_),
    .RESET_B(_00743_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.sum[31] ));
 sky130_fd_sc_hd__dfrtp_1 _11354_ (.CLK(clknet_leaf_100_clk),
    .D(_01919_),
    .RESET_B(_00744_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.sum[32] ));
 sky130_fd_sc_hd__dfrtp_2 _11355_ (.CLK(clknet_leaf_100_clk),
    .D(_01920_),
    .RESET_B(_00745_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.sum[33] ));
 sky130_fd_sc_hd__dfrtp_1 _11356_ (.CLK(clknet_leaf_100_clk),
    .D(_01921_),
    .RESET_B(_00746_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.sum[34] ));
 sky130_fd_sc_hd__dfrtp_1 _11357_ (.CLK(clknet_leaf_100_clk),
    .D(_01922_),
    .RESET_B(_00747_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.sum[35] ));
 sky130_fd_sc_hd__dfrtp_1 _11358_ (.CLK(clknet_leaf_94_clk),
    .D(_01923_),
    .RESET_B(_00748_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.sum[36] ));
 sky130_fd_sc_hd__dfrtp_2 _11359_ (.CLK(clknet_leaf_94_clk),
    .D(_01924_),
    .RESET_B(_00749_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.sum[37] ));
 sky130_fd_sc_hd__dfrtp_2 _11360_ (.CLK(clknet_leaf_94_clk),
    .D(_01925_),
    .RESET_B(_00750_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.sum[38] ));
 sky130_fd_sc_hd__dfrtp_2 _11361_ (.CLK(clknet_leaf_94_clk),
    .D(_01926_),
    .RESET_B(_00751_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.sum[39] ));
 sky130_fd_sc_hd__dfrtp_1 _11362_ (.CLK(clknet_leaf_81_clk),
    .D(_01927_),
    .RESET_B(_00752_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.sum[40] ));
 sky130_fd_sc_hd__dfrtp_2 _11363_ (.CLK(clknet_leaf_91_clk),
    .D(_01928_),
    .RESET_B(_00753_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.sum[41] ));
 sky130_fd_sc_hd__dfrtp_1 _11364_ (.CLK(clknet_leaf_81_clk),
    .D(_01929_),
    .RESET_B(_00754_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.sum[42] ));
 sky130_fd_sc_hd__dfrtp_2 _11365_ (.CLK(clknet_leaf_93_clk),
    .D(_01930_),
    .RESET_B(_00755_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.sum[43] ));
 sky130_fd_sc_hd__dfrtp_2 _11366_ (.CLK(clknet_leaf_93_clk),
    .D(_01931_),
    .RESET_B(_00756_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.sum[44] ));
 sky130_fd_sc_hd__dfrtp_2 _11367_ (.CLK(clknet_leaf_94_clk),
    .D(_01932_),
    .RESET_B(_00757_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.sum[45] ));
 sky130_fd_sc_hd__dfrtp_2 _11368_ (.CLK(clknet_leaf_43_clk),
    .D(_01933_),
    .RESET_B(_00758_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cw1[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11369_ (.CLK(clknet_leaf_41_clk),
    .D(_01934_),
    .RESET_B(_00759_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cw1[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11370_ (.CLK(clknet_leaf_15_clk),
    .D(_01935_),
    .RESET_B(_00760_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cw1[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11371_ (.CLK(clknet_leaf_16_clk),
    .D(_01936_),
    .RESET_B(_00761_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cw1[3] ));
 sky130_fd_sc_hd__dfrtp_2 _11372_ (.CLK(clknet_leaf_15_clk),
    .D(_01937_),
    .RESET_B(_00762_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cw1[4] ));
 sky130_fd_sc_hd__dfrtp_1 _11373_ (.CLK(clknet_leaf_15_clk),
    .D(_01938_),
    .RESET_B(_00763_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cw1[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11374_ (.CLK(clknet_leaf_16_clk),
    .D(_01939_),
    .RESET_B(_00764_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cw1[6] ));
 sky130_fd_sc_hd__dfrtp_1 _11375_ (.CLK(clknet_leaf_13_clk),
    .D(_01940_),
    .RESET_B(_00765_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cw1[7] ));
 sky130_fd_sc_hd__dfrtp_1 _11376_ (.CLK(clknet_leaf_17_clk),
    .D(_01941_),
    .RESET_B(_00766_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cw2[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11377_ (.CLK(clknet_leaf_40_clk),
    .D(_01942_),
    .RESET_B(_00767_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cw2[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11378_ (.CLK(clknet_leaf_17_clk),
    .D(_01943_),
    .RESET_B(_00768_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cw2[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11379_ (.CLK(clknet_leaf_17_clk),
    .D(_01944_),
    .RESET_B(_00769_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cw2[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11380_ (.CLK(clknet_leaf_18_clk),
    .D(_01945_),
    .RESET_B(_00770_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cw2[4] ));
 sky130_fd_sc_hd__dfrtp_1 _11381_ (.CLK(clknet_leaf_19_clk),
    .D(_01946_),
    .RESET_B(_00771_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cw2[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11382_ (.CLK(clknet_leaf_19_clk),
    .D(_01947_),
    .RESET_B(_00772_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cw2[6] ));
 sky130_fd_sc_hd__dfrtp_1 _11383_ (.CLK(clknet_leaf_9_clk),
    .D(_01948_),
    .RESET_B(_00773_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cw2[7] ));
 sky130_fd_sc_hd__dfrtp_4 _11384_ (.CLK(clknet_leaf_15_clk),
    .D(_01949_),
    .RESET_B(_00774_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.histo_index[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11385_ (.CLK(clknet_leaf_15_clk),
    .D(_01950_),
    .RESET_B(_00775_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.histo_index[1] ));
 sky130_fd_sc_hd__dfrtp_4 _11386_ (.CLK(clknet_leaf_15_clk),
    .D(_01951_),
    .RESET_B(_00776_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.histo_index[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11387_ (.CLK(clknet_leaf_15_clk),
    .D(_01952_),
    .RESET_B(_00777_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.histo_index[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11388_ (.CLK(clknet_leaf_15_clk),
    .D(_01953_),
    .RESET_B(_00778_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.histo_index[4] ));
 sky130_fd_sc_hd__dfrtp_1 _11389_ (.CLK(clknet_leaf_14_clk),
    .D(_01954_),
    .RESET_B(_00779_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.histo_index[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11390_ (.CLK(clknet_leaf_14_clk),
    .D(_01955_),
    .RESET_B(_00780_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.histo_index[6] ));
 sky130_fd_sc_hd__dfrtp_4 _11391_ (.CLK(clknet_leaf_13_clk),
    .D(_01956_),
    .RESET_B(_00781_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.histo_index[7] ));
 sky130_fd_sc_hd__dfrtp_4 _11392_ (.CLK(clknet_leaf_13_clk),
    .D(_01957_),
    .RESET_B(_00782_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.histo_index[8] ));
 sky130_fd_sc_hd__dfrtp_1 _11393_ (.CLK(clknet_leaf_12_clk),
    .D(_01958_),
    .RESET_B(_00783_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.controller.fin_FLV ));
 sky130_fd_sc_hd__dfrtp_1 _11394_ (.CLK(clknet_leaf_13_clk),
    .D(_01959_),
    .RESET_B(_00784_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.wipe_the_char_1 ));
 sky130_fd_sc_hd__dfrtp_1 _11395_ (.CLK(clknet_leaf_12_clk),
    .D(_01960_),
    .RESET_B(_00785_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.wipe_the_char_2 ));
 sky130_fd_sc_hd__dfstp_1 _11396_ (.CLK(clknet_leaf_90_clk),
    .D(_01961_),
    .SET_B(_00786_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val1[0] ));
 sky130_fd_sc_hd__dfstp_1 _11397_ (.CLK(clknet_leaf_90_clk),
    .D(_01962_),
    .SET_B(_00787_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val1[1] ));
 sky130_fd_sc_hd__dfstp_1 _11398_ (.CLK(clknet_leaf_90_clk),
    .D(_01963_),
    .SET_B(_00788_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val1[2] ));
 sky130_fd_sc_hd__dfstp_1 _11399_ (.CLK(clknet_leaf_90_clk),
    .D(_01964_),
    .SET_B(_00789_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val1[3] ));
 sky130_fd_sc_hd__dfstp_1 _11400_ (.CLK(clknet_leaf_90_clk),
    .D(_01965_),
    .SET_B(_00790_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val1[4] ));
 sky130_fd_sc_hd__dfstp_1 _11401_ (.CLK(clknet_leaf_91_clk),
    .D(_01966_),
    .SET_B(_00791_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val1[5] ));
 sky130_fd_sc_hd__dfstp_1 _11402_ (.CLK(clknet_leaf_89_clk),
    .D(_01967_),
    .SET_B(_00792_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val1[6] ));
 sky130_fd_sc_hd__dfstp_1 _11403_ (.CLK(clknet_leaf_87_clk),
    .D(_01968_),
    .SET_B(_00793_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val1[7] ));
 sky130_fd_sc_hd__dfstp_2 _11404_ (.CLK(clknet_leaf_87_clk),
    .D(_01969_),
    .SET_B(_00794_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val1[8] ));
 sky130_fd_sc_hd__dfstp_1 _11405_ (.CLK(clknet_leaf_87_clk),
    .D(_01970_),
    .SET_B(_00795_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val1[9] ));
 sky130_fd_sc_hd__dfstp_2 _11406_ (.CLK(clknet_leaf_87_clk),
    .D(_01971_),
    .SET_B(_00796_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val1[10] ));
 sky130_fd_sc_hd__dfstp_1 _11407_ (.CLK(clknet_leaf_87_clk),
    .D(_01972_),
    .SET_B(_00797_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val1[11] ));
 sky130_fd_sc_hd__dfstp_1 _11408_ (.CLK(clknet_leaf_86_clk),
    .D(_01973_),
    .SET_B(_00798_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val1[12] ));
 sky130_fd_sc_hd__dfstp_1 _11409_ (.CLK(clknet_leaf_86_clk),
    .D(_01974_),
    .SET_B(_00799_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val1[13] ));
 sky130_fd_sc_hd__dfstp_1 _11410_ (.CLK(clknet_leaf_85_clk),
    .D(_01975_),
    .SET_B(_00800_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val1[14] ));
 sky130_fd_sc_hd__dfstp_2 _11411_ (.CLK(clknet_leaf_86_clk),
    .D(_01976_),
    .SET_B(_00801_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val1[15] ));
 sky130_fd_sc_hd__dfstp_1 _11412_ (.CLK(clknet_leaf_101_clk),
    .D(_01977_),
    .SET_B(_00802_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val1[16] ));
 sky130_fd_sc_hd__dfstp_2 _11413_ (.CLK(clknet_leaf_101_clk),
    .D(_01978_),
    .SET_B(_00803_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val1[17] ));
 sky130_fd_sc_hd__dfstp_2 _11414_ (.CLK(clknet_leaf_79_clk),
    .D(_01979_),
    .SET_B(_00804_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val1[18] ));
 sky130_fd_sc_hd__dfstp_2 _11415_ (.CLK(clknet_leaf_78_clk),
    .D(_01980_),
    .SET_B(_00805_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val1[19] ));
 sky130_fd_sc_hd__dfstp_1 _11416_ (.CLK(clknet_leaf_78_clk),
    .D(_01981_),
    .SET_B(_00806_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val1[20] ));
 sky130_fd_sc_hd__dfstp_1 _11417_ (.CLK(clknet_leaf_78_clk),
    .D(_01982_),
    .SET_B(_00807_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val1[21] ));
 sky130_fd_sc_hd__dfstp_2 _11418_ (.CLK(clknet_leaf_76_clk),
    .D(_01983_),
    .SET_B(_00808_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val1[22] ));
 sky130_fd_sc_hd__dfstp_2 _11419_ (.CLK(clknet_leaf_76_clk),
    .D(_01984_),
    .SET_B(_00809_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val1[23] ));
 sky130_fd_sc_hd__dfstp_1 _11420_ (.CLK(clknet_leaf_103_clk),
    .D(_01985_),
    .SET_B(_00810_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val1[24] ));
 sky130_fd_sc_hd__dfstp_2 _11421_ (.CLK(clknet_leaf_103_clk),
    .D(_01986_),
    .SET_B(_00811_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val1[25] ));
 sky130_fd_sc_hd__dfstp_2 _11422_ (.CLK(clknet_leaf_103_clk),
    .D(_01987_),
    .SET_B(_00812_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val1[26] ));
 sky130_fd_sc_hd__dfstp_1 _11423_ (.CLK(clknet_leaf_103_clk),
    .D(_01988_),
    .SET_B(_00813_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val1[27] ));
 sky130_fd_sc_hd__dfstp_1 _11424_ (.CLK(clknet_leaf_99_clk),
    .D(_01989_),
    .SET_B(_00814_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val1[28] ));
 sky130_fd_sc_hd__dfstp_2 _11425_ (.CLK(clknet_leaf_99_clk),
    .D(_01990_),
    .SET_B(_00815_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val1[29] ));
 sky130_fd_sc_hd__dfstp_2 _11426_ (.CLK(clknet_leaf_99_clk),
    .D(_01991_),
    .SET_B(_00816_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val1[30] ));
 sky130_fd_sc_hd__dfstp_2 _11427_ (.CLK(clknet_leaf_100_clk),
    .D(_01992_),
    .SET_B(_00817_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val1[31] ));
 sky130_fd_sc_hd__dfstp_1 _11428_ (.CLK(clknet_leaf_98_clk),
    .D(_01993_),
    .SET_B(_00818_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val1[32] ));
 sky130_fd_sc_hd__dfstp_2 _11429_ (.CLK(clknet_leaf_96_clk),
    .D(_01994_),
    .SET_B(_00819_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val1[33] ));
 sky130_fd_sc_hd__dfstp_1 _11430_ (.CLK(clknet_leaf_96_clk),
    .D(_01995_),
    .SET_B(_00820_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val1[34] ));
 sky130_fd_sc_hd__dfstp_2 _11431_ (.CLK(clknet_leaf_96_clk),
    .D(_01996_),
    .SET_B(_00821_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val1[35] ));
 sky130_fd_sc_hd__dfstp_1 _11432_ (.CLK(clknet_leaf_95_clk),
    .D(_01997_),
    .SET_B(_00822_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val1[36] ));
 sky130_fd_sc_hd__dfstp_2 _11433_ (.CLK(clknet_leaf_95_clk),
    .D(_01998_),
    .SET_B(_00823_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val1[37] ));
 sky130_fd_sc_hd__dfstp_2 _11434_ (.CLK(clknet_leaf_95_clk),
    .D(_01999_),
    .SET_B(_00824_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val1[38] ));
 sky130_fd_sc_hd__dfstp_1 _11435_ (.CLK(clknet_leaf_95_clk),
    .D(_02000_),
    .SET_B(_00825_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val1[39] ));
 sky130_fd_sc_hd__dfstp_1 _11436_ (.CLK(clknet_leaf_95_clk),
    .D(_02001_),
    .SET_B(_00826_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val1[40] ));
 sky130_fd_sc_hd__dfstp_1 _11437_ (.CLK(clknet_leaf_95_clk),
    .D(_02002_),
    .SET_B(_00827_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val1[41] ));
 sky130_fd_sc_hd__dfstp_1 _11438_ (.CLK(clknet_leaf_95_clk),
    .D(_02003_),
    .SET_B(_00828_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val1[42] ));
 sky130_fd_sc_hd__dfstp_2 _11439_ (.CLK(clknet_leaf_91_clk),
    .D(_02004_),
    .SET_B(_00829_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val1[43] ));
 sky130_fd_sc_hd__dfstp_1 _11440_ (.CLK(clknet_leaf_93_clk),
    .D(_02005_),
    .SET_B(_00830_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val1[44] ));
 sky130_fd_sc_hd__dfstp_1 _11441_ (.CLK(clknet_leaf_94_clk),
    .D(_02006_),
    .SET_B(_00831_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val1[45] ));
 sky130_fd_sc_hd__dfstp_2 _11442_ (.CLK(clknet_leaf_106_clk),
    .D(_02007_),
    .SET_B(_00832_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val1[46] ));
 sky130_fd_sc_hd__dfstp_1 _11443_ (.CLK(clknet_leaf_90_clk),
    .D(_02008_),
    .SET_B(_00833_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val2[0] ));
 sky130_fd_sc_hd__dfstp_1 _11444_ (.CLK(clknet_leaf_90_clk),
    .D(_02009_),
    .SET_B(_00834_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val2[1] ));
 sky130_fd_sc_hd__dfstp_1 _11445_ (.CLK(clknet_leaf_90_clk),
    .D(_02010_),
    .SET_B(_00835_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val2[2] ));
 sky130_fd_sc_hd__dfstp_1 _11446_ (.CLK(clknet_leaf_89_clk),
    .D(_02011_),
    .SET_B(_00836_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val2[3] ));
 sky130_fd_sc_hd__dfstp_1 _11447_ (.CLK(clknet_leaf_89_clk),
    .D(_02012_),
    .SET_B(_00837_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val2[4] ));
 sky130_fd_sc_hd__dfstp_1 _11448_ (.CLK(clknet_leaf_89_clk),
    .D(_02013_),
    .SET_B(_00838_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val2[5] ));
 sky130_fd_sc_hd__dfstp_1 _11449_ (.CLK(clknet_leaf_88_clk),
    .D(_02014_),
    .SET_B(_00839_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val2[6] ));
 sky130_fd_sc_hd__dfstp_1 _11450_ (.CLK(clknet_leaf_88_clk),
    .D(_02015_),
    .SET_B(_00840_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val2[7] ));
 sky130_fd_sc_hd__dfstp_2 _11451_ (.CLK(clknet_leaf_87_clk),
    .D(_02016_),
    .SET_B(_00841_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val2[8] ));
 sky130_fd_sc_hd__dfstp_1 _11452_ (.CLK(clknet_leaf_88_clk),
    .D(_02017_),
    .SET_B(_00842_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val2[9] ));
 sky130_fd_sc_hd__dfstp_1 _11453_ (.CLK(clknet_leaf_87_clk),
    .D(_02018_),
    .SET_B(_00843_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val2[10] ));
 sky130_fd_sc_hd__dfstp_1 _11454_ (.CLK(clknet_leaf_87_clk),
    .D(_02019_),
    .SET_B(_00844_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val2[11] ));
 sky130_fd_sc_hd__dfstp_1 _11455_ (.CLK(clknet_leaf_86_clk),
    .D(_02020_),
    .SET_B(_00845_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val2[12] ));
 sky130_fd_sc_hd__dfstp_1 _11456_ (.CLK(clknet_leaf_86_clk),
    .D(_02021_),
    .SET_B(_00846_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val2[13] ));
 sky130_fd_sc_hd__dfstp_1 _11457_ (.CLK(clknet_leaf_85_clk),
    .D(_02022_),
    .SET_B(_00847_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val2[14] ));
 sky130_fd_sc_hd__dfstp_2 _11458_ (.CLK(clknet_leaf_79_clk),
    .D(_02023_),
    .SET_B(_00848_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val2[15] ));
 sky130_fd_sc_hd__dfstp_1 _11459_ (.CLK(clknet_leaf_101_clk),
    .D(_02024_),
    .SET_B(_00849_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val2[16] ));
 sky130_fd_sc_hd__dfstp_1 _11460_ (.CLK(clknet_leaf_101_clk),
    .D(_02025_),
    .SET_B(_00850_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val2[17] ));
 sky130_fd_sc_hd__dfstp_2 _11461_ (.CLK(clknet_leaf_79_clk),
    .D(_02026_),
    .SET_B(_00851_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val2[18] ));
 sky130_fd_sc_hd__dfstp_2 _11462_ (.CLK(clknet_leaf_78_clk),
    .D(_02027_),
    .SET_B(_00852_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val2[19] ));
 sky130_fd_sc_hd__dfstp_1 _11463_ (.CLK(clknet_leaf_78_clk),
    .D(_02028_),
    .SET_B(_00853_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val2[20] ));
 sky130_fd_sc_hd__dfstp_1 _11464_ (.CLK(clknet_leaf_78_clk),
    .D(_02029_),
    .SET_B(_00854_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val2[21] ));
 sky130_fd_sc_hd__dfstp_1 _11465_ (.CLK(clknet_leaf_76_clk),
    .D(_02030_),
    .SET_B(_00855_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val2[22] ));
 sky130_fd_sc_hd__dfstp_2 _11466_ (.CLK(clknet_leaf_76_clk),
    .D(_02031_),
    .SET_B(_00856_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val2[23] ));
 sky130_fd_sc_hd__dfstp_2 _11467_ (.CLK(clknet_leaf_102_clk),
    .D(_02032_),
    .SET_B(_00857_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val2[24] ));
 sky130_fd_sc_hd__dfstp_2 _11468_ (.CLK(clknet_leaf_103_clk),
    .D(_02033_),
    .SET_B(_00858_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val2[25] ));
 sky130_fd_sc_hd__dfstp_1 _11469_ (.CLK(clknet_leaf_103_clk),
    .D(_02034_),
    .SET_B(_00859_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val2[26] ));
 sky130_fd_sc_hd__dfstp_1 _11470_ (.CLK(clknet_leaf_102_clk),
    .D(_02035_),
    .SET_B(_00860_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val2[27] ));
 sky130_fd_sc_hd__dfstp_1 _11471_ (.CLK(clknet_leaf_99_clk),
    .D(_02036_),
    .SET_B(_00861_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val2[28] ));
 sky130_fd_sc_hd__dfstp_1 _11472_ (.CLK(clknet_leaf_99_clk),
    .D(_02037_),
    .SET_B(_00862_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val2[29] ));
 sky130_fd_sc_hd__dfstp_2 _11473_ (.CLK(clknet_leaf_99_clk),
    .D(_02038_),
    .SET_B(_00863_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val2[30] ));
 sky130_fd_sc_hd__dfstp_2 _11474_ (.CLK(clknet_leaf_98_clk),
    .D(_02039_),
    .SET_B(_00864_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val2[31] ));
 sky130_fd_sc_hd__dfstp_1 _11475_ (.CLK(clknet_leaf_97_clk),
    .D(_02040_),
    .SET_B(_00865_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val2[32] ));
 sky130_fd_sc_hd__dfstp_1 _11476_ (.CLK(clknet_leaf_97_clk),
    .D(_02041_),
    .SET_B(_00866_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val2[33] ));
 sky130_fd_sc_hd__dfstp_1 _11477_ (.CLK(clknet_leaf_96_clk),
    .D(_02042_),
    .SET_B(_00867_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val2[34] ));
 sky130_fd_sc_hd__dfstp_1 _11478_ (.CLK(clknet_leaf_95_clk),
    .D(_02043_),
    .SET_B(_00868_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val2[35] ));
 sky130_fd_sc_hd__dfstp_1 _11479_ (.CLK(clknet_leaf_95_clk),
    .D(_02044_),
    .SET_B(_00869_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val2[36] ));
 sky130_fd_sc_hd__dfstp_1 _11480_ (.CLK(clknet_leaf_95_clk),
    .D(_02045_),
    .SET_B(_00870_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val2[37] ));
 sky130_fd_sc_hd__dfstp_1 _11481_ (.CLK(clknet_leaf_95_clk),
    .D(_02046_),
    .SET_B(_00871_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val2[38] ));
 sky130_fd_sc_hd__dfstp_1 _11482_ (.CLK(clknet_leaf_95_clk),
    .D(_02047_),
    .SET_B(_00872_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val2[39] ));
 sky130_fd_sc_hd__dfstp_1 _11483_ (.CLK(clknet_leaf_92_clk),
    .D(_02048_),
    .SET_B(_00873_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val2[40] ));
 sky130_fd_sc_hd__dfstp_1 _11484_ (.CLK(clknet_leaf_92_clk),
    .D(_02049_),
    .SET_B(_00874_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val2[41] ));
 sky130_fd_sc_hd__dfstp_1 _11485_ (.CLK(clknet_leaf_91_clk),
    .D(_02050_),
    .SET_B(_00875_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val2[42] ));
 sky130_fd_sc_hd__dfstp_1 _11486_ (.CLK(clknet_leaf_92_clk),
    .D(_02051_),
    .SET_B(_00876_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val2[43] ));
 sky130_fd_sc_hd__dfstp_1 _11487_ (.CLK(clknet_leaf_93_clk),
    .D(_02052_),
    .SET_B(_00877_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val2[44] ));
 sky130_fd_sc_hd__dfstp_1 _11488_ (.CLK(clknet_leaf_94_clk),
    .D(_02053_),
    .SET_B(_00878_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val2[45] ));
 sky130_fd_sc_hd__dfstp_1 _11489_ (.CLK(clknet_leaf_94_clk),
    .D(_02054_),
    .SET_B(_00879_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.val2[46] ));
 sky130_fd_sc_hd__dfstp_1 _11490_ (.CLK(clknet_leaf_12_clk),
    .D(_02055_),
    .SET_B(_00880_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.findLeastValue.startup ));
 sky130_fd_sc_hd__dfrtp_2 _11491_ (.CLK(clknet_leaf_26_clk),
    .D(_02056_),
    .RESET_B(_00881_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.header_synthesis.bit1 ));
 sky130_fd_sc_hd__dfrtp_1 _11492_ (.CLK(clknet_leaf_4_clk),
    .D(_02057_),
    .RESET_B(_00882_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.controller.fin_HG ));
 sky130_fd_sc_hd__dfrtp_1 _11493_ (.CLK(clknet_leaf_3_clk),
    .D(_02058_),
    .RESET_B(_00883_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.total[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11494_ (.CLK(clknet_leaf_2_clk),
    .D(_02059_),
    .RESET_B(_00884_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.total[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11495_ (.CLK(clknet_leaf_0_clk),
    .D(_02060_),
    .RESET_B(_00885_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.total[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11496_ (.CLK(clknet_leaf_119_clk),
    .D(_02061_),
    .RESET_B(_00886_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.total[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11497_ (.CLK(clknet_leaf_119_clk),
    .D(_02062_),
    .RESET_B(_00887_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.total[4] ));
 sky130_fd_sc_hd__dfrtp_1 _11498_ (.CLK(clknet_leaf_0_clk),
    .D(_02063_),
    .RESET_B(_00888_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.total[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11499_ (.CLK(clknet_leaf_0_clk),
    .D(_02064_),
    .RESET_B(_00889_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.total[6] ));
 sky130_fd_sc_hd__dfrtp_1 _11500_ (.CLK(clknet_leaf_120_clk),
    .D(_02065_),
    .RESET_B(_00890_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.total[7] ));
 sky130_fd_sc_hd__dfrtp_1 _11501_ (.CLK(clknet_leaf_120_clk),
    .D(_02066_),
    .RESET_B(_00891_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.total[8] ));
 sky130_fd_sc_hd__dfrtp_1 _11502_ (.CLK(clknet_leaf_120_clk),
    .D(_02067_),
    .RESET_B(_00892_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.total[9] ));
 sky130_fd_sc_hd__dfrtp_1 _11503_ (.CLK(clknet_leaf_120_clk),
    .D(_02068_),
    .RESET_B(_00893_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.total[10] ));
 sky130_fd_sc_hd__dfrtp_1 _11504_ (.CLK(clknet_leaf_120_clk),
    .D(_02069_),
    .RESET_B(_00894_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.total[11] ));
 sky130_fd_sc_hd__dfrtp_1 _11505_ (.CLK(clknet_leaf_119_clk),
    .D(_02070_),
    .RESET_B(_00895_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.total[12] ));
 sky130_fd_sc_hd__dfrtp_1 _11506_ (.CLK(clknet_leaf_118_clk),
    .D(_02071_),
    .RESET_B(_00896_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.total[13] ));
 sky130_fd_sc_hd__dfrtp_1 _11507_ (.CLK(clknet_leaf_119_clk),
    .D(_02072_),
    .RESET_B(_00897_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.total[14] ));
 sky130_fd_sc_hd__dfrtp_1 _11508_ (.CLK(clknet_leaf_119_clk),
    .D(_02073_),
    .RESET_B(_00898_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.total[15] ));
 sky130_fd_sc_hd__dfrtp_1 _11509_ (.CLK(clknet_leaf_119_clk),
    .D(_02074_),
    .RESET_B(_00899_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.total[16] ));
 sky130_fd_sc_hd__dfrtp_1 _11510_ (.CLK(clknet_leaf_119_clk),
    .D(_02075_),
    .RESET_B(_00900_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.total[17] ));
 sky130_fd_sc_hd__dfrtp_1 _11511_ (.CLK(clknet_leaf_117_clk),
    .D(_02076_),
    .RESET_B(_00901_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.total[18] ));
 sky130_fd_sc_hd__dfrtp_1 _11512_ (.CLK(clknet_leaf_118_clk),
    .D(_02077_),
    .RESET_B(_00902_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.total[19] ));
 sky130_fd_sc_hd__dfrtp_1 _11513_ (.CLK(clknet_leaf_117_clk),
    .D(_02078_),
    .RESET_B(_00903_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.total[20] ));
 sky130_fd_sc_hd__dfrtp_1 _11514_ (.CLK(clknet_leaf_118_clk),
    .D(_02079_),
    .RESET_B(_00904_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.total[21] ));
 sky130_fd_sc_hd__dfrtp_1 _11515_ (.CLK(clknet_leaf_118_clk),
    .D(_02080_),
    .RESET_B(_00905_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.total[22] ));
 sky130_fd_sc_hd__dfrtp_1 _11516_ (.CLK(clknet_leaf_118_clk),
    .D(_02081_),
    .RESET_B(_00906_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.total[23] ));
 sky130_fd_sc_hd__dfrtp_1 _11517_ (.CLK(clknet_leaf_118_clk),
    .D(_02082_),
    .RESET_B(_00907_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.total[24] ));
 sky130_fd_sc_hd__dfrtp_1 _11518_ (.CLK(clknet_leaf_119_clk),
    .D(_02083_),
    .RESET_B(_00908_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.total[25] ));
 sky130_fd_sc_hd__dfrtp_1 _11519_ (.CLK(clknet_leaf_119_clk),
    .D(_02084_),
    .RESET_B(_00909_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.total[26] ));
 sky130_fd_sc_hd__dfrtp_1 _11520_ (.CLK(clknet_leaf_119_clk),
    .D(_02085_),
    .RESET_B(_00910_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.total[27] ));
 sky130_fd_sc_hd__dfrtp_1 _11521_ (.CLK(clknet_leaf_119_clk),
    .D(_02086_),
    .RESET_B(_00911_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.total[28] ));
 sky130_fd_sc_hd__dfrtp_1 _11522_ (.CLK(clknet_leaf_120_clk),
    .D(_02087_),
    .RESET_B(_00912_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.total[29] ));
 sky130_fd_sc_hd__dfrtp_1 _11523_ (.CLK(clknet_leaf_120_clk),
    .D(_02088_),
    .RESET_B(_00913_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.total[30] ));
 sky130_fd_sc_hd__dfrtp_1 _11524_ (.CLK(clknet_leaf_120_clk),
    .D(_02089_),
    .RESET_B(_00914_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.total[31] ));
 sky130_fd_sc_hd__dfrtp_1 _11525_ (.CLK(clknet_leaf_80_clk),
    .D(_02090_),
    .RESET_B(_00915_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.sram_out[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11526_ (.CLK(clknet_leaf_80_clk),
    .D(_02091_),
    .RESET_B(_00916_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.sram_out[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11527_ (.CLK(clknet_leaf_80_clk),
    .D(_02092_),
    .RESET_B(_00917_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.sram_out[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11528_ (.CLK(clknet_leaf_85_clk),
    .D(_02093_),
    .RESET_B(_00918_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.sram_out[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11529_ (.CLK(clknet_leaf_81_clk),
    .D(_02094_),
    .RESET_B(_00919_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.sram_out[4] ));
 sky130_fd_sc_hd__dfrtp_1 _11530_ (.CLK(clknet_leaf_81_clk),
    .D(net1465),
    .RESET_B(_00920_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.sram_out[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11531_ (.CLK(clknet_leaf_81_clk),
    .D(_02096_),
    .RESET_B(_00921_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.sram_out[6] ));
 sky130_fd_sc_hd__dfrtp_1 _11532_ (.CLK(clknet_leaf_81_clk),
    .D(_02097_),
    .RESET_B(_00922_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.sram_out[7] ));
 sky130_fd_sc_hd__dfrtp_1 _11533_ (.CLK(clknet_leaf_70_clk),
    .D(_02098_),
    .RESET_B(_00923_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.sram_out[8] ));
 sky130_fd_sc_hd__dfrtp_1 _11534_ (.CLK(clknet_leaf_68_clk),
    .D(_02099_),
    .RESET_B(_00924_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.sram_out[9] ));
 sky130_fd_sc_hd__dfrtp_1 _11535_ (.CLK(clknet_leaf_81_clk),
    .D(_02100_),
    .RESET_B(_00925_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.sram_out[10] ));
 sky130_fd_sc_hd__dfrtp_1 _11536_ (.CLK(clknet_leaf_68_clk),
    .D(_02101_),
    .RESET_B(_00926_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.sram_out[11] ));
 sky130_fd_sc_hd__dfrtp_1 _11537_ (.CLK(clknet_leaf_69_clk),
    .D(_02102_),
    .RESET_B(_00927_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.sram_out[12] ));
 sky130_fd_sc_hd__dfrtp_1 _11538_ (.CLK(clknet_leaf_69_clk),
    .D(_02103_),
    .RESET_B(_00928_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.sram_out[13] ));
 sky130_fd_sc_hd__dfrtp_1 _11539_ (.CLK(clknet_leaf_70_clk),
    .D(_02104_),
    .RESET_B(_00929_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.sram_out[14] ));
 sky130_fd_sc_hd__dfrtp_1 _11540_ (.CLK(clknet_leaf_70_clk),
    .D(_02105_),
    .RESET_B(_00930_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.sram_out[15] ));
 sky130_fd_sc_hd__dfrtp_1 _11541_ (.CLK(clknet_leaf_69_clk),
    .D(_02106_),
    .RESET_B(_00931_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.sram_out[16] ));
 sky130_fd_sc_hd__dfrtp_1 _11542_ (.CLK(clknet_leaf_71_clk),
    .D(_02107_),
    .RESET_B(_00932_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.sram_out[17] ));
 sky130_fd_sc_hd__dfrtp_1 _11543_ (.CLK(clknet_leaf_72_clk),
    .D(_02108_),
    .RESET_B(_00933_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.sram_out[18] ));
 sky130_fd_sc_hd__dfrtp_1 _11544_ (.CLK(clknet_leaf_72_clk),
    .D(_02109_),
    .RESET_B(_00934_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.sram_out[19] ));
 sky130_fd_sc_hd__dfrtp_1 _11545_ (.CLK(clknet_leaf_72_clk),
    .D(_02110_),
    .RESET_B(_00935_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.sram_out[20] ));
 sky130_fd_sc_hd__dfrtp_1 _11546_ (.CLK(clknet_leaf_73_clk),
    .D(_02111_),
    .RESET_B(_00936_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.sram_out[21] ));
 sky130_fd_sc_hd__dfrtp_1 _11547_ (.CLK(clknet_leaf_74_clk),
    .D(_02112_),
    .RESET_B(_00937_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.sram_out[22] ));
 sky130_fd_sc_hd__dfrtp_1 _11548_ (.CLK(clknet_leaf_74_clk),
    .D(_02113_),
    .RESET_B(_00938_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.sram_out[23] ));
 sky130_fd_sc_hd__dfrtp_1 _11549_ (.CLK(clknet_leaf_47_clk),
    .D(_02114_),
    .RESET_B(_00939_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.sram_out[24] ));
 sky130_fd_sc_hd__dfrtp_1 _11550_ (.CLK(clknet_leaf_45_clk),
    .D(_02115_),
    .RESET_B(_00940_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.sram_out[25] ));
 sky130_fd_sc_hd__dfrtp_1 _11551_ (.CLK(clknet_leaf_46_clk),
    .D(_02116_),
    .RESET_B(_00941_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.sram_out[26] ));
 sky130_fd_sc_hd__dfrtp_1 _11552_ (.CLK(clknet_leaf_46_clk),
    .D(_02117_),
    .RESET_B(_00942_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.sram_out[27] ));
 sky130_fd_sc_hd__dfrtp_1 _11553_ (.CLK(clknet_leaf_42_clk),
    .D(_02118_),
    .RESET_B(_00943_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.sram_out[28] ));
 sky130_fd_sc_hd__dfrtp_1 _11554_ (.CLK(clknet_leaf_41_clk),
    .D(_02119_),
    .RESET_B(_00944_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.sram_out[29] ));
 sky130_fd_sc_hd__dfrtp_1 _11555_ (.CLK(clknet_leaf_41_clk),
    .D(_02120_),
    .RESET_B(_00945_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.sram_out[30] ));
 sky130_fd_sc_hd__dfrtp_1 _11556_ (.CLK(clknet_leaf_40_clk),
    .D(_02121_),
    .RESET_B(_00946_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.sram_out[31] ));
 sky130_fd_sc_hd__dfrtp_1 _11557_ (.CLK(clknet_leaf_7_clk),
    .D(_02122_),
    .RESET_B(_00947_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net64));
 sky130_fd_sc_hd__dfrtp_1 _11558_ (.CLK(clknet_leaf_21_clk),
    .D(_02123_),
    .RESET_B(_00948_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net65));
 sky130_fd_sc_hd__dfrtp_1 _11559_ (.CLK(clknet_leaf_21_clk),
    .D(_02124_),
    .RESET_B(_00949_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net66));
 sky130_fd_sc_hd__dfrtp_1 _11560_ (.CLK(clknet_leaf_21_clk),
    .D(_02125_),
    .RESET_B(_00950_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net67));
 sky130_fd_sc_hd__dfrtp_2 _11561_ (.CLK(clknet_leaf_21_clk),
    .D(_02126_),
    .RESET_B(_00951_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net68));
 sky130_fd_sc_hd__dfrtp_1 _11562_ (.CLK(clknet_leaf_21_clk),
    .D(_02127_),
    .RESET_B(_00952_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net69));
 sky130_fd_sc_hd__dfrtp_1 _11563_ (.CLK(clknet_leaf_6_clk),
    .D(_02128_),
    .RESET_B(_00953_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net70));
 sky130_fd_sc_hd__dfrtp_1 _11564_ (.CLK(clknet_leaf_6_clk),
    .D(_02129_),
    .RESET_B(_00954_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net71));
 sky130_fd_sc_hd__dfrtp_1 _11565_ (.CLK(clknet_leaf_7_clk),
    .D(_02130_),
    .RESET_B(_00955_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net45));
 sky130_fd_sc_hd__dfrtp_1 _11566_ (.CLK(clknet_leaf_5_clk),
    .D(_02131_),
    .RESET_B(_00956_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net46));
 sky130_fd_sc_hd__dfrtp_1 _11567_ (.CLK(clknet_leaf_6_clk),
    .D(_02132_),
    .RESET_B(_00957_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net47));
 sky130_fd_sc_hd__dfrtp_1 _11568_ (.CLK(clknet_leaf_7_clk),
    .D(_02133_),
    .RESET_B(_00958_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net48));
 sky130_fd_sc_hd__dfrtp_1 _11569_ (.CLK(clknet_leaf_23_clk),
    .D(_02134_),
    .RESET_B(_00959_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net49));
 sky130_fd_sc_hd__dfrtp_1 _11570_ (.CLK(clknet_leaf_27_clk),
    .D(_02135_),
    .RESET_B(_00960_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net50));
 sky130_fd_sc_hd__dfrtp_1 _11571_ (.CLK(clknet_leaf_27_clk),
    .D(_02136_),
    .RESET_B(_00961_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net51));
 sky130_fd_sc_hd__dfrtp_1 _11572_ (.CLK(clknet_leaf_5_clk),
    .D(_02137_),
    .RESET_B(_00962_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net52));
 sky130_fd_sc_hd__dfrtp_1 _11573_ (.CLK(clknet_leaf_31_clk),
    .D(_02138_),
    .RESET_B(_00963_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net53));
 sky130_fd_sc_hd__dfrtp_1 _11574_ (.CLK(clknet_leaf_27_clk),
    .D(_02139_),
    .RESET_B(_00964_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net54));
 sky130_fd_sc_hd__dfrtp_1 _11575_ (.CLK(clknet_leaf_31_clk),
    .D(_02140_),
    .RESET_B(_00965_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net55));
 sky130_fd_sc_hd__dfrtp_1 _11576_ (.CLK(clknet_leaf_27_clk),
    .D(_02141_),
    .RESET_B(_00966_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net56));
 sky130_fd_sc_hd__dfrtp_1 _11577_ (.CLK(clknet_leaf_27_clk),
    .D(_02142_),
    .RESET_B(_00967_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net57));
 sky130_fd_sc_hd__dfrtp_1 _11578_ (.CLK(clknet_leaf_5_clk),
    .D(_02143_),
    .RESET_B(_00968_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net58));
 sky130_fd_sc_hd__dfrtp_1 _11579_ (.CLK(clknet_leaf_6_clk),
    .D(_02144_),
    .RESET_B(_00969_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net59));
 sky130_fd_sc_hd__dfrtp_1 _11580_ (.CLK(clknet_leaf_5_clk),
    .D(_02145_),
    .RESET_B(_00970_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net60));
 sky130_fd_sc_hd__dfrtp_1 _11581_ (.CLK(clknet_leaf_27_clk),
    .D(_02146_),
    .RESET_B(_00971_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net61));
 sky130_fd_sc_hd__dfrtp_1 _11582_ (.CLK(clknet_leaf_5_clk),
    .D(_02147_),
    .RESET_B(_00972_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net63));
 sky130_fd_sc_hd__dfrtp_1 _11583_ (.CLK(clknet_leaf_4_clk),
    .D(_02148_),
    .RESET_B(_00973_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.out_of_init ));
 sky130_fd_sc_hd__dfrtp_1 _11584_ (.CLK(clknet_leaf_30_clk),
    .D(_02149_),
    .RESET_B(_00974_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.count[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11585_ (.CLK(clknet_leaf_30_clk),
    .D(_02150_),
    .RESET_B(_00975_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11586_ (.CLK(clknet_leaf_30_clk),
    .D(_02151_),
    .RESET_B(_00976_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11587_ (.CLK(clknet_leaf_30_clk),
    .D(_02152_),
    .RESET_B(_00977_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.count[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11588_ (.CLK(clknet_leaf_31_clk),
    .D(_02153_),
    .RESET_B(_00978_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.count[4] ));
 sky130_fd_sc_hd__dfrtp_1 _11589_ (.CLK(clknet_leaf_30_clk),
    .D(_02154_),
    .RESET_B(_00979_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.count[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11590_ (.CLK(clknet_leaf_32_clk),
    .D(_02155_),
    .RESET_B(_00980_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.count[6] ));
 sky130_fd_sc_hd__dfrtp_1 _11591_ (.CLK(clknet_leaf_31_clk),
    .D(_02156_),
    .RESET_B(_00981_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.cb_syn.count[7] ));
 sky130_fd_sc_hd__dfrtp_1 _11592_ (.CLK(clknet_leaf_4_clk),
    .D(\top.dut.out_valid_next ),
    .RESET_B(_00982_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.dut.out_valid ));
 sky130_fd_sc_hd__dfrtp_1 _11593_ (.CLK(clknet_leaf_0_clk),
    .D(\top.dut.bit_buf_next[0] ),
    .RESET_B(_00983_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.dut.bit_buf[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11594_ (.CLK(clknet_leaf_5_clk),
    .D(\top.dut.bit_buf_next[1] ),
    .RESET_B(_00984_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.dut.bit_buf[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11595_ (.CLK(clknet_leaf_0_clk),
    .D(\top.dut.bit_buf_next[2] ),
    .RESET_B(_00985_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.dut.bit_buf[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11596_ (.CLK(clknet_leaf_5_clk),
    .D(\top.dut.bit_buf_next[3] ),
    .RESET_B(_00986_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.dut.bit_buf[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11597_ (.CLK(clknet_leaf_120_clk),
    .D(\top.dut.bit_buf_next[4] ),
    .RESET_B(_00987_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.dut.bit_buf[4] ));
 sky130_fd_sc_hd__dfrtp_1 _11598_ (.CLK(clknet_leaf_120_clk),
    .D(\top.dut.bit_buf_next[5] ),
    .RESET_B(_00988_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.dut.bit_buf[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11599_ (.CLK(clknet_leaf_0_clk),
    .D(\top.dut.bit_buf_next[6] ),
    .RESET_B(_00989_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.dut.bit_buf[6] ));
 sky130_fd_sc_hd__dfrtp_1 _11600_ (.CLK(clknet_leaf_0_clk),
    .D(\top.dut.bit_buf_next[7] ),
    .RESET_B(_00990_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.dut.bit_buf[7] ));
 sky130_fd_sc_hd__dfrtp_1 _11601_ (.CLK(clknet_leaf_1_clk),
    .D(\top.dut.bit_buf_next[8] ),
    .RESET_B(_00991_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.dut.bit_buf[8] ));
 sky130_fd_sc_hd__dfrtp_1 _11602_ (.CLK(clknet_leaf_0_clk),
    .D(\top.dut.bit_buf_next[9] ),
    .RESET_B(_00992_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.dut.bit_buf[9] ));
 sky130_fd_sc_hd__dfrtp_1 _11603_ (.CLK(clknet_leaf_5_clk),
    .D(\top.dut.bit_buf_next[10] ),
    .RESET_B(_00993_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.dut.bit_buf[10] ));
 sky130_fd_sc_hd__dfrtp_1 _11604_ (.CLK(clknet_leaf_120_clk),
    .D(\top.dut.bit_buf_next[11] ),
    .RESET_B(_00994_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.dut.bit_buf[11] ));
 sky130_fd_sc_hd__dfrtp_1 _11605_ (.CLK(clknet_leaf_120_clk),
    .D(\top.dut.bit_buf_next[12] ),
    .RESET_B(_00995_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.dut.bit_buf[12] ));
 sky130_fd_sc_hd__dfrtp_1 _11606_ (.CLK(clknet_leaf_0_clk),
    .D(\top.dut.bit_buf_next[13] ),
    .RESET_B(_00996_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.dut.bit_buf[13] ));
 sky130_fd_sc_hd__dfrtp_1 _11607_ (.CLK(clknet_leaf_7_clk),
    .D(_02157_),
    .RESET_B(_00997_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.sram_interface.check ));
 sky130_fd_sc_hd__dfrtp_4 _11608_ (.CLK(clknet_leaf_22_clk),
    .D(_02158_),
    .RESET_B(_00998_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.sram_interface.init_counter[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11609_ (.CLK(clknet_leaf_21_clk),
    .D(_02159_),
    .RESET_B(_00999_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.sram_interface.init_counter[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11610_ (.CLK(clknet_leaf_22_clk),
    .D(_02160_),
    .RESET_B(_01000_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.sram_interface.init_counter[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11611_ (.CLK(clknet_leaf_22_clk),
    .D(_02161_),
    .RESET_B(_01001_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.sram_interface.init_counter[3] ));
 sky130_fd_sc_hd__dfrtp_2 _11612_ (.CLK(clknet_leaf_22_clk),
    .D(_02162_),
    .RESET_B(_01002_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.sram_interface.init_counter[4] ));
 sky130_fd_sc_hd__dfrtp_1 _11613_ (.CLK(clknet_leaf_22_clk),
    .D(_02163_),
    .RESET_B(_01003_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.sram_interface.init_counter[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11614_ (.CLK(clknet_leaf_22_clk),
    .D(_02164_),
    .RESET_B(_01004_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.sram_interface.init_counter[6] ));
 sky130_fd_sc_hd__dfrtp_4 _11615_ (.CLK(clknet_leaf_22_clk),
    .D(_02165_),
    .RESET_B(_01005_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.sram_interface.init_counter[7] ));
 sky130_fd_sc_hd__dfrtp_1 _11616_ (.CLK(clknet_leaf_24_clk),
    .D(_02166_),
    .RESET_B(_01006_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.sram_interface.init_counter[8] ));
 sky130_fd_sc_hd__dfrtp_1 _11617_ (.CLK(clknet_leaf_22_clk),
    .D(_02167_),
    .RESET_B(_01007_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.sram_interface.init_counter[9] ));
 sky130_fd_sc_hd__dfrtp_2 _11618_ (.CLK(clknet_leaf_22_clk),
    .D(_02168_),
    .RESET_B(_01008_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.sram_interface.init_counter[10] ));
 sky130_fd_sc_hd__dfrtp_1 _11619_ (.CLK(clknet_leaf_22_clk),
    .D(net1102),
    .RESET_B(_01009_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.sram_interface.init_counter[11] ));
 sky130_fd_sc_hd__dfrtp_1 _11620_ (.CLK(clknet_leaf_28_clk),
    .D(_02170_),
    .RESET_B(_01010_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.sram_interface.init_counter[12] ));
 sky130_fd_sc_hd__dfrtp_1 _11621_ (.CLK(clknet_leaf_28_clk),
    .D(_02171_),
    .RESET_B(_01011_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.sram_interface.init_counter[13] ));
 sky130_fd_sc_hd__dfrtp_1 _11622_ (.CLK(clknet_leaf_28_clk),
    .D(_02172_),
    .RESET_B(_01012_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.sram_interface.init_counter[14] ));
 sky130_fd_sc_hd__dfrtp_1 _11623_ (.CLK(clknet_leaf_28_clk),
    .D(_02173_),
    .RESET_B(_01013_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.sram_interface.init_counter[15] ));
 sky130_fd_sc_hd__dfrtp_1 _11624_ (.CLK(clknet_leaf_23_clk),
    .D(_02174_),
    .RESET_B(_01014_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.sram_interface.init_counter[16] ));
 sky130_fd_sc_hd__dfrtp_1 _11625_ (.CLK(clknet_leaf_23_clk),
    .D(_02175_),
    .RESET_B(_01015_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.sram_interface.init_counter[17] ));
 sky130_fd_sc_hd__dfrtp_1 _11626_ (.CLK(clknet_leaf_23_clk),
    .D(_02176_),
    .RESET_B(_01016_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.sram_interface.init_counter[18] ));
 sky130_fd_sc_hd__dfrtp_1 _11627_ (.CLK(clknet_leaf_23_clk),
    .D(_02177_),
    .RESET_B(_01017_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.sram_interface.init_counter[19] ));
 sky130_fd_sc_hd__dfrtp_1 _11628_ (.CLK(clknet_leaf_28_clk),
    .D(_02178_),
    .RESET_B(_01018_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.sram_interface.init_counter[20] ));
 sky130_fd_sc_hd__dfrtp_1 _11629_ (.CLK(clknet_leaf_28_clk),
    .D(_02179_),
    .RESET_B(_01019_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.sram_interface.init_counter[21] ));
 sky130_fd_sc_hd__dfrtp_1 _11630_ (.CLK(clknet_leaf_29_clk),
    .D(_02180_),
    .RESET_B(_01020_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.sram_interface.init_counter[22] ));
 sky130_fd_sc_hd__dfrtp_1 _11631_ (.CLK(clknet_leaf_28_clk),
    .D(_02181_),
    .RESET_B(_01021_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.sram_interface.init_counter[23] ));
 sky130_fd_sc_hd__dfrtp_1 _11632_ (.CLK(clknet_leaf_10_clk),
    .D(_02182_),
    .RESET_B(_01022_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.TRN_sram_complete ));
 sky130_fd_sc_hd__dfrtp_1 _11633_ (.CLK(clknet_leaf_110_clk),
    .D(_02183_),
    .RESET_B(_01023_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[32] ));
 sky130_fd_sc_hd__dfrtp_1 _11634_ (.CLK(clknet_leaf_110_clk),
    .D(_02184_),
    .RESET_B(_01024_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[33] ));
 sky130_fd_sc_hd__dfrtp_1 _11635_ (.CLK(clknet_leaf_98_clk),
    .D(_02185_),
    .RESET_B(_01025_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[34] ));
 sky130_fd_sc_hd__dfrtp_1 _11636_ (.CLK(clknet_leaf_97_clk),
    .D(_02186_),
    .RESET_B(_01026_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[35] ));
 sky130_fd_sc_hd__dfrtp_1 _11637_ (.CLK(clknet_leaf_98_clk),
    .D(_02187_),
    .RESET_B(_01027_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[36] ));
 sky130_fd_sc_hd__dfrtp_1 _11638_ (.CLK(clknet_leaf_100_clk),
    .D(_02188_),
    .RESET_B(_01028_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[37] ));
 sky130_fd_sc_hd__dfrtp_1 _11639_ (.CLK(clknet_leaf_98_clk),
    .D(_02189_),
    .RESET_B(_01029_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[38] ));
 sky130_fd_sc_hd__dfrtp_1 _11640_ (.CLK(clknet_leaf_110_clk),
    .D(_02190_),
    .RESET_B(_01030_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[39] ));
 sky130_fd_sc_hd__dfrtp_1 _11641_ (.CLK(clknet_leaf_109_clk),
    .D(_02191_),
    .RESET_B(_01031_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[40] ));
 sky130_fd_sc_hd__dfrtp_1 _11642_ (.CLK(clknet_leaf_110_clk),
    .D(_02192_),
    .RESET_B(_01032_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[41] ));
 sky130_fd_sc_hd__dfrtp_1 _11643_ (.CLK(clknet_leaf_109_clk),
    .D(_02193_),
    .RESET_B(_01033_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[42] ));
 sky130_fd_sc_hd__dfrtp_1 _11644_ (.CLK(clknet_leaf_109_clk),
    .D(_02194_),
    .RESET_B(_01034_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[43] ));
 sky130_fd_sc_hd__dfrtp_1 _11645_ (.CLK(clknet_leaf_109_clk),
    .D(_02195_),
    .RESET_B(_01035_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[44] ));
 sky130_fd_sc_hd__dfrtp_1 _11646_ (.CLK(clknet_leaf_108_clk),
    .D(_02196_),
    .RESET_B(_01036_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[45] ));
 sky130_fd_sc_hd__dfrtp_1 _11647_ (.CLK(clknet_leaf_111_clk),
    .D(_02197_),
    .RESET_B(_01037_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[46] ));
 sky130_fd_sc_hd__dfrtp_1 _11648_ (.CLK(clknet_leaf_111_clk),
    .D(_02198_),
    .RESET_B(_01038_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[47] ));
 sky130_fd_sc_hd__dfrtp_1 _11649_ (.CLK(clknet_leaf_115_clk),
    .D(_02199_),
    .RESET_B(_01039_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[48] ));
 sky130_fd_sc_hd__dfrtp_1 _11650_ (.CLK(clknet_leaf_115_clk),
    .D(_02200_),
    .RESET_B(_01040_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[49] ));
 sky130_fd_sc_hd__dfrtp_1 _11651_ (.CLK(clknet_leaf_115_clk),
    .D(_02201_),
    .RESET_B(_01041_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[50] ));
 sky130_fd_sc_hd__dfrtp_1 _11652_ (.CLK(clknet_leaf_115_clk),
    .D(_02202_),
    .RESET_B(_01042_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[51] ));
 sky130_fd_sc_hd__dfrtp_1 _11653_ (.CLK(clknet_leaf_115_clk),
    .D(_02203_),
    .RESET_B(_01043_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[52] ));
 sky130_fd_sc_hd__dfrtp_1 _11654_ (.CLK(clknet_leaf_115_clk),
    .D(_02204_),
    .RESET_B(_01044_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[53] ));
 sky130_fd_sc_hd__dfrtp_1 _11655_ (.CLK(clknet_leaf_114_clk),
    .D(_02205_),
    .RESET_B(_01045_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[54] ));
 sky130_fd_sc_hd__dfrtp_1 _11656_ (.CLK(clknet_leaf_115_clk),
    .D(_02206_),
    .RESET_B(_01046_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[55] ));
 sky130_fd_sc_hd__dfrtp_1 _11657_ (.CLK(clknet_leaf_114_clk),
    .D(_02207_),
    .RESET_B(_01047_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[56] ));
 sky130_fd_sc_hd__dfrtp_1 _11658_ (.CLK(clknet_leaf_114_clk),
    .D(_02208_),
    .RESET_B(_01048_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[57] ));
 sky130_fd_sc_hd__dfrtp_1 _11659_ (.CLK(clknet_leaf_117_clk),
    .D(_02209_),
    .RESET_B(_01049_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[58] ));
 sky130_fd_sc_hd__dfrtp_1 _11660_ (.CLK(clknet_leaf_114_clk),
    .D(_02210_),
    .RESET_B(_01050_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[59] ));
 sky130_fd_sc_hd__dfrtp_1 _11661_ (.CLK(clknet_leaf_115_clk),
    .D(_02211_),
    .RESET_B(_01051_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[60] ));
 sky130_fd_sc_hd__dfrtp_1 _11662_ (.CLK(clknet_leaf_114_clk),
    .D(_02212_),
    .RESET_B(_01052_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[61] ));
 sky130_fd_sc_hd__dfrtp_1 _11663_ (.CLK(clknet_leaf_113_clk),
    .D(_02213_),
    .RESET_B(_01053_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[62] ));
 sky130_fd_sc_hd__dfrtp_1 _11664_ (.CLK(clknet_leaf_113_clk),
    .D(_02214_),
    .RESET_B(_01054_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.path[63] ));
 sky130_fd_sc_hd__dfrtp_4 _11665_ (.CLK(clknet_leaf_19_clk),
    .D(_02215_),
    .RESET_B(_01055_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.CB_write_complete ));
 sky130_fd_sc_hd__dfrtp_2 _11666_ (.CLK(clknet_leaf_18_clk),
    .D(_02216_),
    .RESET_B(_01056_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.CB_read_complete ));
 sky130_fd_sc_hd__dfrtp_2 _11667_ (.CLK(clknet_leaf_91_clk),
    .D(_02217_),
    .RESET_B(_01057_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.compVal[0] ));
 sky130_fd_sc_hd__dfrtp_2 _11668_ (.CLK(clknet_leaf_91_clk),
    .D(_02218_),
    .RESET_B(_01058_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.compVal[1] ));
 sky130_fd_sc_hd__dfrtp_2 _11669_ (.CLK(clknet_leaf_91_clk),
    .D(_02219_),
    .RESET_B(_01059_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.compVal[2] ));
 sky130_fd_sc_hd__dfrtp_2 _11670_ (.CLK(clknet_leaf_91_clk),
    .D(_02220_),
    .RESET_B(_01060_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.compVal[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11671_ (.CLK(clknet_leaf_91_clk),
    .D(_02221_),
    .RESET_B(_01061_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.compVal[4] ));
 sky130_fd_sc_hd__dfrtp_2 _11672_ (.CLK(clknet_leaf_93_clk),
    .D(_02222_),
    .RESET_B(_01062_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.compVal[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11673_ (.CLK(clknet_leaf_93_clk),
    .D(_02223_),
    .RESET_B(_01063_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.compVal[6] ));
 sky130_fd_sc_hd__dfrtp_1 _11674_ (.CLK(clknet_leaf_93_clk),
    .D(_02224_),
    .RESET_B(_01064_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.compVal[7] ));
 sky130_fd_sc_hd__dfrtp_2 _11675_ (.CLK(clknet_leaf_87_clk),
    .D(_02225_),
    .RESET_B(_01065_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.compVal[8] ));
 sky130_fd_sc_hd__dfrtp_2 _11676_ (.CLK(clknet_leaf_87_clk),
    .D(_02226_),
    .RESET_B(_01066_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.compVal[9] ));
 sky130_fd_sc_hd__dfrtp_4 _11677_ (.CLK(clknet_leaf_91_clk),
    .D(_02227_),
    .RESET_B(_01067_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.compVal[10] ));
 sky130_fd_sc_hd__dfrtp_1 _11678_ (.CLK(clknet_leaf_86_clk),
    .D(_02228_),
    .RESET_B(_01068_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.compVal[11] ));
 sky130_fd_sc_hd__dfrtp_2 _11679_ (.CLK(clknet_leaf_86_clk),
    .D(_02229_),
    .RESET_B(_01069_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.compVal[12] ));
 sky130_fd_sc_hd__dfrtp_2 _11680_ (.CLK(clknet_leaf_94_clk),
    .D(_02230_),
    .RESET_B(_01070_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.compVal[13] ));
 sky130_fd_sc_hd__dfrtp_4 _11681_ (.CLK(clknet_leaf_86_clk),
    .D(_02231_),
    .RESET_B(_01071_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.compVal[14] ));
 sky130_fd_sc_hd__dfrtp_1 _11682_ (.CLK(clknet_leaf_94_clk),
    .D(_02232_),
    .RESET_B(_01072_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.compVal[15] ));
 sky130_fd_sc_hd__dfrtp_2 _11683_ (.CLK(clknet_leaf_100_clk),
    .D(_02233_),
    .RESET_B(_01073_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.compVal[16] ));
 sky130_fd_sc_hd__dfrtp_1 _11684_ (.CLK(clknet_leaf_94_clk),
    .D(_02234_),
    .RESET_B(_01074_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.compVal[17] ));
 sky130_fd_sc_hd__dfrtp_4 _11685_ (.CLK(clknet_leaf_100_clk),
    .D(_02235_),
    .RESET_B(_01075_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.compVal[18] ));
 sky130_fd_sc_hd__dfrtp_4 _11686_ (.CLK(clknet_leaf_100_clk),
    .D(_02236_),
    .RESET_B(_01076_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.compVal[19] ));
 sky130_fd_sc_hd__dfrtp_4 _11687_ (.CLK(clknet_leaf_102_clk),
    .D(_02237_),
    .RESET_B(_01077_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.compVal[20] ));
 sky130_fd_sc_hd__dfrtp_2 _11688_ (.CLK(clknet_leaf_78_clk),
    .D(_02238_),
    .RESET_B(_01078_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.compVal[21] ));
 sky130_fd_sc_hd__dfrtp_2 _11689_ (.CLK(clknet_leaf_76_clk),
    .D(_02239_),
    .RESET_B(_01079_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.compVal[22] ));
 sky130_fd_sc_hd__dfrtp_2 _11690_ (.CLK(clknet_leaf_76_clk),
    .D(_02240_),
    .RESET_B(_01080_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.compVal[23] ));
 sky130_fd_sc_hd__dfrtp_2 _11691_ (.CLK(clknet_leaf_102_clk),
    .D(_02241_),
    .RESET_B(_01081_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.compVal[24] ));
 sky130_fd_sc_hd__dfrtp_2 _11692_ (.CLK(clknet_leaf_103_clk),
    .D(_02242_),
    .RESET_B(_01082_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.compVal[25] ));
 sky130_fd_sc_hd__dfrtp_4 _11693_ (.CLK(clknet_leaf_103_clk),
    .D(_02243_),
    .RESET_B(_01083_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.compVal[26] ));
 sky130_fd_sc_hd__dfrtp_2 _11694_ (.CLK(clknet_leaf_103_clk),
    .D(_02244_),
    .RESET_B(_01084_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.compVal[27] ));
 sky130_fd_sc_hd__dfrtp_2 _11695_ (.CLK(clknet_leaf_99_clk),
    .D(_02245_),
    .RESET_B(_01085_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.compVal[28] ));
 sky130_fd_sc_hd__dfrtp_2 _11696_ (.CLK(clknet_leaf_98_clk),
    .D(_02246_),
    .RESET_B(_01086_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.compVal[29] ));
 sky130_fd_sc_hd__dfrtp_1 _11697_ (.CLK(clknet_leaf_110_clk),
    .D(_02247_),
    .RESET_B(_01087_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.compVal[30] ));
 sky130_fd_sc_hd__dfrtp_1 _11698_ (.CLK(clknet_leaf_98_clk),
    .D(_02248_),
    .RESET_B(_01088_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.compVal[31] ));
 sky130_fd_sc_hd__dfrtp_2 _11699_ (.CLK(clknet_leaf_9_clk),
    .D(_02249_),
    .RESET_B(_01089_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.sram_interface.CB_write_counter[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11700_ (.CLK(clknet_leaf_8_clk),
    .D(_02250_),
    .RESET_B(_01090_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.sram_interface.CB_write_counter[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11701_ (.CLK(clknet_leaf_19_clk),
    .D(net957),
    .RESET_B(_01091_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.sram_interface.CB_read_counter ));
 sky130_fd_sc_hd__dfrtp_2 _11702_ (.CLK(clknet_leaf_85_clk),
    .D(_02252_),
    .RESET_B(_01092_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hist_data_o[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11703_ (.CLK(clknet_leaf_80_clk),
    .D(_02253_),
    .RESET_B(_01093_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hist_data_o[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11704_ (.CLK(clknet_leaf_80_clk),
    .D(_02254_),
    .RESET_B(_01094_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hist_data_o[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11705_ (.CLK(clknet_leaf_80_clk),
    .D(_02255_),
    .RESET_B(_01095_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hist_data_o[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11706_ (.CLK(clknet_leaf_80_clk),
    .D(_02256_),
    .RESET_B(_01096_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hist_data_o[4] ));
 sky130_fd_sc_hd__dfrtp_1 _11707_ (.CLK(clknet_leaf_80_clk),
    .D(_02257_),
    .RESET_B(_01097_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hist_data_o[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11708_ (.CLK(clknet_leaf_80_clk),
    .D(_02258_),
    .RESET_B(_01098_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hist_data_o[6] ));
 sky130_fd_sc_hd__dfrtp_1 _11709_ (.CLK(clknet_leaf_80_clk),
    .D(_02259_),
    .RESET_B(_01099_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hist_data_o[7] ));
 sky130_fd_sc_hd__dfrtp_1 _11710_ (.CLK(clknet_leaf_81_clk),
    .D(_02260_),
    .RESET_B(_01100_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hist_data_o[8] ));
 sky130_fd_sc_hd__dfrtp_1 _11711_ (.CLK(clknet_leaf_81_clk),
    .D(_02261_),
    .RESET_B(_01101_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hist_data_o[9] ));
 sky130_fd_sc_hd__dfrtp_1 _11712_ (.CLK(clknet_leaf_81_clk),
    .D(_02262_),
    .RESET_B(_01102_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hist_data_o[10] ));
 sky130_fd_sc_hd__dfrtp_1 _11713_ (.CLK(clknet_leaf_69_clk),
    .D(_02263_),
    .RESET_B(_01103_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hist_data_o[11] ));
 sky130_fd_sc_hd__dfrtp_1 _11714_ (.CLK(clknet_leaf_69_clk),
    .D(_02264_),
    .RESET_B(_01104_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hist_data_o[12] ));
 sky130_fd_sc_hd__dfrtp_1 _11715_ (.CLK(clknet_leaf_69_clk),
    .D(_02265_),
    .RESET_B(_01105_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hist_data_o[13] ));
 sky130_fd_sc_hd__dfrtp_1 _11716_ (.CLK(clknet_leaf_69_clk),
    .D(_02266_),
    .RESET_B(_01106_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hist_data_o[14] ));
 sky130_fd_sc_hd__dfrtp_1 _11717_ (.CLK(clknet_leaf_70_clk),
    .D(_02267_),
    .RESET_B(_01107_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hist_data_o[15] ));
 sky130_fd_sc_hd__dfrtp_1 _11718_ (.CLK(clknet_leaf_73_clk),
    .D(_02268_),
    .RESET_B(_01108_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hist_data_o[16] ));
 sky130_fd_sc_hd__dfrtp_1 _11719_ (.CLK(clknet_leaf_73_clk),
    .D(_02269_),
    .RESET_B(_01109_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hist_data_o[17] ));
 sky130_fd_sc_hd__dfrtp_1 _11720_ (.CLK(clknet_leaf_72_clk),
    .D(_02270_),
    .RESET_B(_01110_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hist_data_o[18] ));
 sky130_fd_sc_hd__dfrtp_1 _11721_ (.CLK(clknet_leaf_72_clk),
    .D(_02271_),
    .RESET_B(_01111_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hist_data_o[19] ));
 sky130_fd_sc_hd__dfrtp_1 _11722_ (.CLK(clknet_leaf_72_clk),
    .D(_02272_),
    .RESET_B(_01112_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hist_data_o[20] ));
 sky130_fd_sc_hd__dfrtp_1 _11723_ (.CLK(clknet_leaf_74_clk),
    .D(_02273_),
    .RESET_B(_01113_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hist_data_o[21] ));
 sky130_fd_sc_hd__dfrtp_1 _11724_ (.CLK(clknet_leaf_74_clk),
    .D(_02274_),
    .RESET_B(_01114_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hist_data_o[22] ));
 sky130_fd_sc_hd__dfrtp_1 _11725_ (.CLK(clknet_leaf_45_clk),
    .D(_02275_),
    .RESET_B(_01115_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hist_data_o[23] ));
 sky130_fd_sc_hd__dfrtp_1 _11726_ (.CLK(clknet_leaf_47_clk),
    .D(_02276_),
    .RESET_B(_01116_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hist_data_o[24] ));
 sky130_fd_sc_hd__dfrtp_1 _11727_ (.CLK(clknet_leaf_45_clk),
    .D(_02277_),
    .RESET_B(_01117_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hist_data_o[25] ));
 sky130_fd_sc_hd__dfrtp_1 _11728_ (.CLK(clknet_leaf_46_clk),
    .D(_02278_),
    .RESET_B(_01118_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hist_data_o[26] ));
 sky130_fd_sc_hd__dfrtp_1 _11729_ (.CLK(clknet_leaf_42_clk),
    .D(_02279_),
    .RESET_B(_01119_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hist_data_o[27] ));
 sky130_fd_sc_hd__dfrtp_1 _11730_ (.CLK(clknet_leaf_41_clk),
    .D(_02280_),
    .RESET_B(_01120_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hist_data_o[28] ));
 sky130_fd_sc_hd__dfrtp_1 _11731_ (.CLK(clknet_leaf_40_clk),
    .D(_02281_),
    .RESET_B(_01121_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hist_data_o[29] ));
 sky130_fd_sc_hd__dfrtp_1 _11732_ (.CLK(clknet_leaf_40_clk),
    .D(_02282_),
    .RESET_B(_01122_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hist_data_o[30] ));
 sky130_fd_sc_hd__dfrtp_1 _11733_ (.CLK(clknet_leaf_40_clk),
    .D(_02283_),
    .RESET_B(_01123_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hist_data_o[31] ));
 sky130_fd_sc_hd__dfrtp_4 _11734_ (.CLK(clknet_leaf_12_clk),
    .D(_02284_),
    .RESET_B(_01124_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.write_HT_fin ));
 sky130_fd_sc_hd__dfrtp_1 _11735_ (.CLK(clknet_leaf_12_clk),
    .D(_02285_),
    .RESET_B(_01125_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.FLV_done ));
 sky130_fd_sc_hd__dfstp_1 _11736_ (.CLK(clknet_leaf_7_clk),
    .D(_02286_),
    .SET_B(_01126_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.init ));
 sky130_fd_sc_hd__dfrtp_1 _11737_ (.CLK(clknet_leaf_107_clk),
    .D(_02287_),
    .RESET_B(_01127_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.sram_interface.counter_HTREE[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11738_ (.CLK(clknet_leaf_106_clk),
    .D(_02288_),
    .RESET_B(_01128_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.sram_interface.counter_HTREE[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11739_ (.CLK(clknet_leaf_107_clk),
    .D(_02289_),
    .RESET_B(_01129_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.sram_interface.counter_HTREE[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11740_ (.CLK(clknet_leaf_106_clk),
    .D(_02290_),
    .RESET_B(_01130_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.sram_interface.counter_HTREE[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11741_ (.CLK(clknet_leaf_4_clk),
    .D(_02291_),
    .RESET_B(_01131_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.sram_interface.write_counter_FLV[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11742_ (.CLK(clknet_leaf_4_clk),
    .D(_02292_),
    .RESET_B(_01132_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.sram_interface.write_counter_FLV[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11743_ (.CLK(clknet_leaf_10_clk),
    .D(_02293_),
    .RESET_B(_01133_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.sram_interface.write_counter_FLV[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11744_ (.CLK(clknet_leaf_6_clk),
    .D(_02294_),
    .RESET_B(_01134_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.histogram.init_edge ));
 sky130_fd_sc_hd__dfrtp_1 _11745_ (.CLK(clknet_leaf_11_clk),
    .D(_02295_),
    .RESET_B(_01135_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.sram_interface.zero_cnt[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11746_ (.CLK(clknet_leaf_11_clk),
    .D(_02296_),
    .RESET_B(_01136_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.sram_interface.zero_cnt[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11747_ (.CLK(clknet_leaf_11_clk),
    .D(_02297_),
    .RESET_B(_01137_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.sram_interface.zero_cnt[2] ));
 sky130_fd_sc_hd__dfstp_1 _11748_ (.CLK(clknet_leaf_106_clk),
    .D(_00017_),
    .SET_B(_01138_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11749_ (.CLK(clknet_leaf_106_clk),
    .D(_00019_),
    .RESET_B(_01139_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11750_ (.CLK(clknet_leaf_105_clk),
    .D(net1638),
    .RESET_B(_01140_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.state[2] ));
 sky130_fd_sc_hd__dfrtp_2 _11751_ (.CLK(clknet_leaf_104_clk),
    .D(_00021_),
    .RESET_B(_01141_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.state[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11752_ (.CLK(clknet_leaf_105_clk),
    .D(_00022_),
    .RESET_B(_01142_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.state[4] ));
 sky130_fd_sc_hd__dfrtp_1 _11753_ (.CLK(clknet_leaf_105_clk),
    .D(net1523),
    .RESET_B(_01143_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.state[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11754_ (.CLK(clknet_leaf_105_clk),
    .D(_00024_),
    .RESET_B(_01144_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.state[6] ));
 sky130_fd_sc_hd__dfrtp_1 _11755_ (.CLK(clknet_leaf_105_clk),
    .D(_00025_),
    .RESET_B(_01145_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.state[7] ));
 sky130_fd_sc_hd__dfrtp_1 _11756_ (.CLK(clknet_leaf_105_clk),
    .D(_00026_),
    .RESET_B(_01146_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.state[8] ));
 sky130_fd_sc_hd__dfrtp_1 _11757_ (.CLK(clknet_leaf_105_clk),
    .D(net1543),
    .RESET_B(_01147_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.state[9] ));
 sky130_fd_sc_hd__dfrtp_1 _11758_ (.CLK(clknet_leaf_106_clk),
    .D(_00018_),
    .RESET_B(_01148_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.state[10] ));
 sky130_fd_sc_hd__dfxtp_1 _11759_ (.CLK(clknet_leaf_47_clk),
    .D(_02298_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[46] ));
 sky130_fd_sc_hd__dfxtp_1 _11760_ (.CLK(clknet_leaf_46_clk),
    .D(_02299_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[47] ));
 sky130_fd_sc_hd__dfxtp_1 _11761_ (.CLK(clknet_leaf_45_clk),
    .D(_02300_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[48] ));
 sky130_fd_sc_hd__dfxtp_1 _11762_ (.CLK(clknet_leaf_74_clk),
    .D(net1276),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[49] ));
 sky130_fd_sc_hd__dfxtp_1 _11763_ (.CLK(clknet_leaf_72_clk),
    .D(_02302_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[50] ));
 sky130_fd_sc_hd__dfxtp_1 _11764_ (.CLK(clknet_leaf_47_clk),
    .D(_02303_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[51] ));
 sky130_fd_sc_hd__dfxtp_1 _11765_ (.CLK(clknet_leaf_72_clk),
    .D(_02304_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[52] ));
 sky130_fd_sc_hd__dfxtp_1 _11766_ (.CLK(clknet_leaf_72_clk),
    .D(_02305_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[53] ));
 sky130_fd_sc_hd__dfxtp_1 _11767_ (.CLK(clknet_leaf_76_clk),
    .D(_02306_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[54] ));
 sky130_fd_sc_hd__dfxtp_1 _11768_ (.CLK(clknet_leaf_74_clk),
    .D(_02307_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[55] ));
 sky130_fd_sc_hd__dfxtp_1 _11769_ (.CLK(clknet_leaf_45_clk),
    .D(_02308_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[56] ));
 sky130_fd_sc_hd__dfxtp_1 _11770_ (.CLK(clknet_leaf_45_clk),
    .D(_02309_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[57] ));
 sky130_fd_sc_hd__dfxtp_1 _11771_ (.CLK(clknet_leaf_74_clk),
    .D(net991),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[58] ));
 sky130_fd_sc_hd__dfxtp_1 _11772_ (.CLK(clknet_leaf_75_clk),
    .D(_02311_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[59] ));
 sky130_fd_sc_hd__dfxtp_1 _11773_ (.CLK(clknet_leaf_42_clk),
    .D(_02312_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[60] ));
 sky130_fd_sc_hd__dfxtp_1 _11774_ (.CLK(clknet_leaf_41_clk),
    .D(_02313_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[61] ));
 sky130_fd_sc_hd__dfxtp_1 _11775_ (.CLK(clknet_leaf_41_clk),
    .D(_02314_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[62] ));
 sky130_fd_sc_hd__dfxtp_1 _11776_ (.CLK(clknet_leaf_75_clk),
    .D(_02315_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.hTree.node_reg[63] ));
 sky130_fd_sc_hd__dfrtp_4 _11777_ (.CLK(clknet_leaf_3_clk),
    .D(_00012_),
    .RESET_B(_01149_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.controller.state_reg[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11778_ (.CLK(clknet_leaf_3_clk),
    .D(_00013_),
    .RESET_B(_01150_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.controller.state_reg[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11779_ (.CLK(clknet_leaf_3_clk),
    .D(_00014_),
    .RESET_B(_01151_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.controller.state_reg[4] ));
 sky130_fd_sc_hd__dfrtp_2 _11780_ (.CLK(clknet_leaf_3_clk),
    .D(_00015_),
    .RESET_B(_01152_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.controller.state_reg[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11781_ (.CLK(clknet_leaf_3_clk),
    .D(_00016_),
    .RESET_B(_01153_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.sram_interface.write_HT_fin_n ));
 sky130_fd_sc_hd__dfrtp_1 _11782_ (.CLK(clknet_leaf_2_clk),
    .D(_02316_),
    .RESET_B(_01154_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.translation.write_fin ));
 sky130_fd_sc_hd__dfrtp_4 _11783_ (.CLK(clknet_leaf_97_clk),
    .D(_02317_),
    .RESET_B(_01155_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.compVal[32] ));
 sky130_fd_sc_hd__dfrtp_2 _11784_ (.CLK(clknet_leaf_96_clk),
    .D(_02318_),
    .RESET_B(_01156_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.compVal[33] ));
 sky130_fd_sc_hd__dfrtp_2 _11785_ (.CLK(clknet_leaf_96_clk),
    .D(_02319_),
    .RESET_B(_01157_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.compVal[34] ));
 sky130_fd_sc_hd__dfrtp_4 _11786_ (.CLK(clknet_leaf_96_clk),
    .D(_02320_),
    .RESET_B(_01158_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.compVal[35] ));
 sky130_fd_sc_hd__dfrtp_2 _11787_ (.CLK(clknet_leaf_95_clk),
    .D(_02321_),
    .RESET_B(_01159_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.compVal[36] ));
 sky130_fd_sc_hd__dfrtp_4 _11788_ (.CLK(clknet_leaf_95_clk),
    .D(_02322_),
    .RESET_B(_01160_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.compVal[37] ));
 sky130_fd_sc_hd__dfrtp_2 _11789_ (.CLK(clknet_leaf_95_clk),
    .D(_02323_),
    .RESET_B(_01161_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.compVal[38] ));
 sky130_fd_sc_hd__dfrtp_2 _11790_ (.CLK(clknet_leaf_95_clk),
    .D(_02324_),
    .RESET_B(_01162_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.compVal[39] ));
 sky130_fd_sc_hd__dfrtp_4 _11791_ (.CLK(clknet_leaf_92_clk),
    .D(_02325_),
    .RESET_B(_01163_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.compVal[40] ));
 sky130_fd_sc_hd__dfrtp_4 _11792_ (.CLK(clknet_leaf_92_clk),
    .D(_02326_),
    .RESET_B(_01164_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.compVal[41] ));
 sky130_fd_sc_hd__dfrtp_2 _11793_ (.CLK(clknet_leaf_92_clk),
    .D(_02327_),
    .RESET_B(_01165_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.compVal[42] ));
 sky130_fd_sc_hd__dfrtp_1 _11794_ (.CLK(clknet_leaf_92_clk),
    .D(_02328_),
    .RESET_B(_01166_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.compVal[43] ));
 sky130_fd_sc_hd__dfrtp_2 _11795_ (.CLK(clknet_leaf_92_clk),
    .D(_02329_),
    .RESET_B(_01167_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.compVal[44] ));
 sky130_fd_sc_hd__dfrtp_2 _11796_ (.CLK(clknet_leaf_94_clk),
    .D(_02330_),
    .RESET_B(_01168_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.compVal[45] ));
 sky130_fd_sc_hd__dfrtp_4 _11797_ (.CLK(clknet_leaf_119_clk),
    .D(net441),
    .RESET_B(_01169_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.WB.prev_BUSY_O ));
 sky130_fd_sc_hd__dfrtp_4 _11798_ (.CLK(clknet_leaf_5_clk),
    .D(_02331_),
    .RESET_B(_01170_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.TRN_char_index[0] ));
 sky130_fd_sc_hd__dfrtp_4 _11799_ (.CLK(clknet_leaf_7_clk),
    .D(_02332_),
    .RESET_B(_01171_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.TRN_char_index[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11800_ (.CLK(clknet_leaf_6_clk),
    .D(_02333_),
    .RESET_B(_01172_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.TRN_char_index[2] ));
 sky130_fd_sc_hd__dfrtp_2 _11801_ (.CLK(clknet_leaf_7_clk),
    .D(_02334_),
    .RESET_B(_01173_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.TRN_char_index[3] ));
 sky130_fd_sc_hd__dfrtp_4 _11802_ (.CLK(clknet_leaf_6_clk),
    .D(_02335_),
    .RESET_B(_01174_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.TRN_char_index[4] ));
 sky130_fd_sc_hd__dfrtp_4 _11803_ (.CLK(clknet_leaf_5_clk),
    .D(_02336_),
    .RESET_B(_01175_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.TRN_char_index[5] ));
 sky130_fd_sc_hd__dfrtp_4 _11804_ (.CLK(clknet_leaf_4_clk),
    .D(_02337_),
    .RESET_B(_01176_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.TRN_char_index[6] ));
 sky130_fd_sc_hd__dfrtp_1 _11805_ (.CLK(clknet_leaf_83_clk),
    .D(_02338_),
    .RESET_B(_01177_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net73));
 sky130_fd_sc_hd__dfrtp_1 _11806_ (.CLK(clknet_leaf_83_clk),
    .D(_02339_),
    .RESET_B(_01178_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net84));
 sky130_fd_sc_hd__dfrtp_1 _11807_ (.CLK(clknet_leaf_83_clk),
    .D(_02340_),
    .RESET_B(_01179_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net95));
 sky130_fd_sc_hd__dfrtp_1 _11808_ (.CLK(clknet_leaf_83_clk),
    .D(_02341_),
    .RESET_B(_01180_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net98));
 sky130_fd_sc_hd__dfrtp_1 _11809_ (.CLK(clknet_leaf_83_clk),
    .D(_02342_),
    .RESET_B(_01181_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net99));
 sky130_fd_sc_hd__dfrtp_1 _11810_ (.CLK(clknet_leaf_82_clk),
    .D(_02343_),
    .RESET_B(_01182_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net100));
 sky130_fd_sc_hd__dfrtp_1 _11811_ (.CLK(clknet_leaf_82_clk),
    .D(_02344_),
    .RESET_B(_01183_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net101));
 sky130_fd_sc_hd__dfrtp_1 _11812_ (.CLK(clknet_leaf_82_clk),
    .D(_02345_),
    .RESET_B(_01184_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net102));
 sky130_fd_sc_hd__dfrtp_1 _11813_ (.CLK(clknet_leaf_65_clk),
    .D(_02346_),
    .RESET_B(_01185_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net103));
 sky130_fd_sc_hd__dfrtp_1 _11814_ (.CLK(clknet_leaf_82_clk),
    .D(_02347_),
    .RESET_B(_01186_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net104));
 sky130_fd_sc_hd__dfrtp_1 _11815_ (.CLK(clknet_leaf_67_clk),
    .D(_02348_),
    .RESET_B(_01187_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net74));
 sky130_fd_sc_hd__dfrtp_1 _11816_ (.CLK(clknet_leaf_67_clk),
    .D(_02349_),
    .RESET_B(_01188_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net75));
 sky130_fd_sc_hd__dfrtp_1 _11817_ (.CLK(clknet_leaf_66_clk),
    .D(_02350_),
    .RESET_B(_01189_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net76));
 sky130_fd_sc_hd__dfrtp_1 _11818_ (.CLK(clknet_leaf_66_clk),
    .D(_02351_),
    .RESET_B(_01190_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net77));
 sky130_fd_sc_hd__dfrtp_1 _11819_ (.CLK(clknet_leaf_65_clk),
    .D(_02352_),
    .RESET_B(_01191_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net78));
 sky130_fd_sc_hd__dfrtp_1 _11820_ (.CLK(clknet_leaf_65_clk),
    .D(_02353_),
    .RESET_B(_01192_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net79));
 sky130_fd_sc_hd__dfrtp_1 _11821_ (.CLK(clknet_leaf_66_clk),
    .D(_02354_),
    .RESET_B(_01193_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net80));
 sky130_fd_sc_hd__dfrtp_1 _11822_ (.CLK(clknet_leaf_66_clk),
    .D(_02355_),
    .RESET_B(_01194_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net81));
 sky130_fd_sc_hd__dfrtp_1 _11823_ (.CLK(clknet_leaf_65_clk),
    .D(_02356_),
    .RESET_B(_01195_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net82));
 sky130_fd_sc_hd__dfrtp_1 _11824_ (.CLK(clknet_leaf_65_clk),
    .D(_02357_),
    .RESET_B(_01196_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net83));
 sky130_fd_sc_hd__dfrtp_1 _11825_ (.CLK(clknet_leaf_66_clk),
    .D(_02358_),
    .RESET_B(_01197_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net85));
 sky130_fd_sc_hd__dfrtp_1 _11826_ (.CLK(clknet_leaf_65_clk),
    .D(_02359_),
    .RESET_B(_01198_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net86));
 sky130_fd_sc_hd__dfrtp_1 _11827_ (.CLK(clknet_leaf_66_clk),
    .D(_02360_),
    .RESET_B(_01199_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net87));
 sky130_fd_sc_hd__dfrtp_1 _11828_ (.CLK(clknet_leaf_67_clk),
    .D(_02361_),
    .RESET_B(_01200_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net88));
 sky130_fd_sc_hd__dfrtp_1 _11829_ (.CLK(clknet_leaf_47_clk),
    .D(_02362_),
    .RESET_B(_01201_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net89));
 sky130_fd_sc_hd__dfrtp_1 _11830_ (.CLK(clknet_leaf_67_clk),
    .D(_02363_),
    .RESET_B(_01202_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net90));
 sky130_fd_sc_hd__dfrtp_1 _11831_ (.CLK(clknet_leaf_67_clk),
    .D(_02364_),
    .RESET_B(_01203_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net91));
 sky130_fd_sc_hd__dfrtp_1 _11832_ (.CLK(clknet_leaf_82_clk),
    .D(_02365_),
    .RESET_B(_01204_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net92));
 sky130_fd_sc_hd__dfrtp_1 _11833_ (.CLK(clknet_leaf_46_clk),
    .D(_02366_),
    .RESET_B(_01205_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net93));
 sky130_fd_sc_hd__dfrtp_1 _11834_ (.CLK(clknet_leaf_42_clk),
    .D(_02367_),
    .RESET_B(_01206_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net94));
 sky130_fd_sc_hd__dfrtp_1 _11835_ (.CLK(clknet_leaf_41_clk),
    .D(_02368_),
    .RESET_B(_01207_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net96));
 sky130_fd_sc_hd__dfrtp_1 _11836_ (.CLK(clknet_leaf_41_clk),
    .D(_02369_),
    .RESET_B(_01208_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net97));
 sky130_fd_sc_hd__dfrtp_2 _11837_ (.CLK(clknet_leaf_5_clk),
    .D(_02370_),
    .RESET_B(_01209_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net72));
 sky130_fd_sc_hd__dfrtp_1 _11838_ (.CLK(clknet_leaf_65_clk),
    .D(_02371_),
    .RESET_B(_01210_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net110));
 sky130_fd_sc_hd__dfrtp_4 _11839_ (.CLK(clknet_leaf_96_clk),
    .D(_02372_),
    .RESET_B(_01211_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.WB.CPU_DAT_O[0] ));
 sky130_fd_sc_hd__dfrtp_4 _11840_ (.CLK(clknet_leaf_113_clk),
    .D(_02373_),
    .RESET_B(_01212_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.WB.CPU_DAT_O[1] ));
 sky130_fd_sc_hd__dfrtp_4 _11841_ (.CLK(clknet_leaf_112_clk),
    .D(_02374_),
    .RESET_B(_01213_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.WB.CPU_DAT_O[2] ));
 sky130_fd_sc_hd__dfrtp_4 _11842_ (.CLK(clknet_leaf_112_clk),
    .D(_02375_),
    .RESET_B(_01214_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.WB.CPU_DAT_O[3] ));
 sky130_fd_sc_hd__dfrtp_4 _11843_ (.CLK(clknet_leaf_96_clk),
    .D(_02376_),
    .RESET_B(_01215_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.WB.CPU_DAT_O[4] ));
 sky130_fd_sc_hd__dfrtp_4 _11844_ (.CLK(clknet_leaf_113_clk),
    .D(_02377_),
    .RESET_B(_01216_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.WB.CPU_DAT_O[5] ));
 sky130_fd_sc_hd__dfrtp_4 _11845_ (.CLK(clknet_leaf_96_clk),
    .D(_02378_),
    .RESET_B(_01217_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.WB.CPU_DAT_O[6] ));
 sky130_fd_sc_hd__dfrtp_4 _11846_ (.CLK(clknet_leaf_96_clk),
    .D(_02379_),
    .RESET_B(_01218_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.WB.CPU_DAT_O[7] ));
 sky130_fd_sc_hd__dfrtp_4 _11847_ (.CLK(clknet_leaf_114_clk),
    .D(_02380_),
    .RESET_B(_01219_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.WB.CPU_DAT_O[8] ));
 sky130_fd_sc_hd__dfrtp_4 _11848_ (.CLK(clknet_leaf_112_clk),
    .D(_02381_),
    .RESET_B(_01220_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.WB.CPU_DAT_O[9] ));
 sky130_fd_sc_hd__dfrtp_4 _11849_ (.CLK(clknet_leaf_114_clk),
    .D(_02382_),
    .RESET_B(_01221_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.WB.CPU_DAT_O[10] ));
 sky130_fd_sc_hd__dfrtp_4 _11850_ (.CLK(clknet_leaf_96_clk),
    .D(_02383_),
    .RESET_B(_01222_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.WB.CPU_DAT_O[11] ));
 sky130_fd_sc_hd__dfrtp_4 _11851_ (.CLK(clknet_leaf_96_clk),
    .D(_02384_),
    .RESET_B(_01223_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.WB.CPU_DAT_O[12] ));
 sky130_fd_sc_hd__dfrtp_4 _11852_ (.CLK(clknet_leaf_112_clk),
    .D(_02385_),
    .RESET_B(_01224_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.WB.CPU_DAT_O[13] ));
 sky130_fd_sc_hd__dfrtp_4 _11853_ (.CLK(clknet_leaf_114_clk),
    .D(_02386_),
    .RESET_B(_01225_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.WB.CPU_DAT_O[14] ));
 sky130_fd_sc_hd__dfrtp_4 _11854_ (.CLK(clknet_leaf_97_clk),
    .D(_02387_),
    .RESET_B(_01226_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.WB.CPU_DAT_O[15] ));
 sky130_fd_sc_hd__dfrtp_4 _11855_ (.CLK(clknet_leaf_96_clk),
    .D(_02388_),
    .RESET_B(_01227_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.WB.CPU_DAT_O[16] ));
 sky130_fd_sc_hd__dfrtp_4 _11856_ (.CLK(clknet_leaf_112_clk),
    .D(_02389_),
    .RESET_B(_01228_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.WB.CPU_DAT_O[17] ));
 sky130_fd_sc_hd__dfrtp_4 _11857_ (.CLK(clknet_leaf_112_clk),
    .D(_02390_),
    .RESET_B(_01229_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.WB.CPU_DAT_O[18] ));
 sky130_fd_sc_hd__dfrtp_4 _11858_ (.CLK(clknet_leaf_113_clk),
    .D(_02391_),
    .RESET_B(_01230_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.WB.CPU_DAT_O[19] ));
 sky130_fd_sc_hd__dfrtp_4 _11859_ (.CLK(clknet_leaf_96_clk),
    .D(_02392_),
    .RESET_B(_01231_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.WB.CPU_DAT_O[20] ));
 sky130_fd_sc_hd__dfrtp_4 _11860_ (.CLK(clknet_leaf_114_clk),
    .D(_02393_),
    .RESET_B(_01232_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.WB.CPU_DAT_O[21] ));
 sky130_fd_sc_hd__dfrtp_4 _11861_ (.CLK(clknet_leaf_112_clk),
    .D(_02394_),
    .RESET_B(_01233_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.WB.CPU_DAT_O[22] ));
 sky130_fd_sc_hd__dfrtp_4 _11862_ (.CLK(clknet_leaf_112_clk),
    .D(_02395_),
    .RESET_B(_01234_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.WB.CPU_DAT_O[23] ));
 sky130_fd_sc_hd__dfrtp_4 _11863_ (.CLK(clknet_leaf_113_clk),
    .D(_02396_),
    .RESET_B(_01235_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.WB.CPU_DAT_O[24] ));
 sky130_fd_sc_hd__dfrtp_4 _11864_ (.CLK(clknet_leaf_113_clk),
    .D(_02397_),
    .RESET_B(_01236_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.WB.CPU_DAT_O[25] ));
 sky130_fd_sc_hd__dfrtp_4 _11865_ (.CLK(clknet_leaf_113_clk),
    .D(_02398_),
    .RESET_B(_01237_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.WB.CPU_DAT_O[26] ));
 sky130_fd_sc_hd__dfrtp_4 _11866_ (.CLK(clknet_leaf_112_clk),
    .D(_02399_),
    .RESET_B(_01238_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.WB.CPU_DAT_O[27] ));
 sky130_fd_sc_hd__dfrtp_4 _11867_ (.CLK(clknet_leaf_112_clk),
    .D(_02400_),
    .RESET_B(_01239_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.WB.CPU_DAT_O[28] ));
 sky130_fd_sc_hd__dfrtp_4 _11868_ (.CLK(clknet_leaf_112_clk),
    .D(_02401_),
    .RESET_B(_01240_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.WB.CPU_DAT_O[29] ));
 sky130_fd_sc_hd__dfrtp_4 _11869_ (.CLK(clknet_leaf_113_clk),
    .D(_02402_),
    .RESET_B(_01241_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.WB.CPU_DAT_O[30] ));
 sky130_fd_sc_hd__dfrtp_4 _11870_ (.CLK(clknet_leaf_112_clk),
    .D(_02403_),
    .RESET_B(_01242_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.WB.CPU_DAT_O[31] ));
 sky130_fd_sc_hd__dfrtp_4 _11871_ (.CLK(clknet_leaf_26_clk),
    .D(\top.header_synthesis.next_write_num_lefts ),
    .RESET_B(_01243_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.header_synthesis.write_num_lefts ));
 sky130_fd_sc_hd__dfrtp_1 _11872_ (.CLK(clknet_leaf_1_clk),
    .D(\top.dut.bits_in_buf_next[0] ),
    .RESET_B(_01244_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.dut.bits_in_buf[0] ));
 sky130_fd_sc_hd__dfrtp_2 _11873_ (.CLK(clknet_leaf_1_clk),
    .D(\top.dut.bits_in_buf_next[1] ),
    .RESET_B(_01245_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.dut.bits_in_buf[1] ));
 sky130_fd_sc_hd__dfrtp_4 _11874_ (.CLK(clknet_leaf_1_clk),
    .D(\top.dut.bits_in_buf_next[2] ),
    .RESET_B(_01246_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.dut.bits_in_buf[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11875_ (.CLK(clknet_leaf_120_clk),
    .D(net878),
    .RESET_B(_01247_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\top.dut.bits_in_buf[3] ));
 sky130_fd_sc_hd__buf_2 _11876_ (.A(net879),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ADR_O[0]));
 sky130_fd_sc_hd__buf_2 _11877_ (.A(net880),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ADR_O[1]));
 sky130_fd_sc_hd__buf_2 _11878_ (.A(net881),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ADR_O[27]));
 sky130_fd_sc_hd__clkbuf_1 _11879_ (.A(net63),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net62));
 sky130_fd_sc_hd__buf_2 _11880_ (.A(net882),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ADR_O[30]));
 sky130_fd_sc_hd__buf_2 _11881_ (.A(net883),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ADR_O[31]));
 sky130_fd_sc_hd__clkbuf_1 _11882_ (.A(net441),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_1 _11883_ (.A(net441),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_1 _11884_ (.A(net441),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_1 _11885_ (.A(net441),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_1 _11886_ (.A(net441),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net109));
 sky130_fd_sc_hd__buf_2 _11887_ (.A(net919),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_oeb[0]));
 sky130_fd_sc_hd__buf_2 _11888_ (.A(net884),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_oeb[1]));
 sky130_fd_sc_hd__buf_2 _11889_ (.A(net920),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_oeb[2]));
 sky130_fd_sc_hd__buf_2 _11890_ (.A(net921),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_oeb[3]));
 sky130_fd_sc_hd__buf_2 _11891_ (.A(net922),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_oeb[4]));
 sky130_fd_sc_hd__buf_2 _11892_ (.A(net923),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_oeb[5]));
 sky130_fd_sc_hd__buf_2 _11893_ (.A(net924),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_oeb[6]));
 sky130_fd_sc_hd__buf_2 _11894_ (.A(net925),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_oeb[7]));
 sky130_fd_sc_hd__buf_2 _11895_ (.A(net926),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_oeb[8]));
 sky130_fd_sc_hd__buf_2 _11896_ (.A(net927),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_oeb[9]));
 sky130_fd_sc_hd__buf_2 _11897_ (.A(net928),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_oeb[10]));
 sky130_fd_sc_hd__buf_2 _11898_ (.A(net929),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_oeb[11]));
 sky130_fd_sc_hd__buf_2 _11899_ (.A(net930),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_oeb[12]));
 sky130_fd_sc_hd__buf_2 _11900_ (.A(net931),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_oeb[13]));
 sky130_fd_sc_hd__buf_2 _11901_ (.A(net932),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_oeb[14]));
 sky130_fd_sc_hd__buf_2 _11902_ (.A(net933),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_oeb[15]));
 sky130_fd_sc_hd__buf_2 _11903_ (.A(net934),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_oeb[16]));
 sky130_fd_sc_hd__buf_2 _11904_ (.A(net935),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_oeb[17]));
 sky130_fd_sc_hd__buf_2 _11905_ (.A(net936),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_oeb[18]));
 sky130_fd_sc_hd__buf_2 _11906_ (.A(net937),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_oeb[19]));
 sky130_fd_sc_hd__buf_2 _11907_ (.A(net938),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_oeb[20]));
 sky130_fd_sc_hd__buf_2 _11908_ (.A(net939),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_oeb[21]));
 sky130_fd_sc_hd__buf_2 _11909_ (.A(net940),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_oeb[22]));
 sky130_fd_sc_hd__buf_2 _11910_ (.A(net941),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_oeb[23]));
 sky130_fd_sc_hd__buf_2 _11911_ (.A(net942),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_oeb[24]));
 sky130_fd_sc_hd__buf_2 _11912_ (.A(net943),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_oeb[25]));
 sky130_fd_sc_hd__buf_2 _11913_ (.A(net944),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_oeb[26]));
 sky130_fd_sc_hd__buf_2 _11914_ (.A(net945),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_oeb[27]));
 sky130_fd_sc_hd__buf_2 _11915_ (.A(net946),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_oeb[28]));
 sky130_fd_sc_hd__buf_2 _11916_ (.A(net947),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_oeb[29]));
 sky130_fd_sc_hd__buf_2 _11917_ (.A(net948),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_oeb[30]));
 sky130_fd_sc_hd__buf_2 _11918_ (.A(net949),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_oeb[31]));
 sky130_fd_sc_hd__buf_2 _11919_ (.A(net950),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_oeb[32]));
 sky130_fd_sc_hd__buf_2 _11920_ (.A(net951),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_oeb[33]));
 sky130_fd_sc_hd__buf_2 _11921_ (.A(net885),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_out[0]));
 sky130_fd_sc_hd__clkbuf_1 _11922_ (.A(\top.translation.writeBin ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net111));
 sky130_fd_sc_hd__buf_2 _11923_ (.A(net886),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_out[2]));
 sky130_fd_sc_hd__buf_2 _11924_ (.A(net887),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_out[3]));
 sky130_fd_sc_hd__buf_2 _11925_ (.A(net888),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_out[4]));
 sky130_fd_sc_hd__buf_2 _11926_ (.A(net889),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_out[5]));
 sky130_fd_sc_hd__buf_2 _11927_ (.A(net890),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_out[6]));
 sky130_fd_sc_hd__buf_2 _11928_ (.A(net891),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_out[7]));
 sky130_fd_sc_hd__buf_2 _11929_ (.A(net892),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_out[8]));
 sky130_fd_sc_hd__buf_2 _11930_ (.A(net893),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_out[9]));
 sky130_fd_sc_hd__buf_2 _11931_ (.A(net894),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_out[10]));
 sky130_fd_sc_hd__buf_2 _11932_ (.A(net895),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_out[11]));
 sky130_fd_sc_hd__buf_2 _11933_ (.A(net896),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_out[12]));
 sky130_fd_sc_hd__buf_2 _11934_ (.A(net897),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_out[13]));
 sky130_fd_sc_hd__buf_2 _11935_ (.A(net898),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_out[14]));
 sky130_fd_sc_hd__buf_2 _11936_ (.A(net899),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_out[15]));
 sky130_fd_sc_hd__buf_2 _11937_ (.A(net900),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_out[16]));
 sky130_fd_sc_hd__buf_2 _11938_ (.A(net901),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_out[17]));
 sky130_fd_sc_hd__buf_2 _11939_ (.A(net902),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_out[18]));
 sky130_fd_sc_hd__buf_2 _11940_ (.A(net903),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_out[19]));
 sky130_fd_sc_hd__buf_2 _11941_ (.A(net904),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_out[20]));
 sky130_fd_sc_hd__buf_2 _11942_ (.A(net905),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_out[21]));
 sky130_fd_sc_hd__buf_2 _11943_ (.A(net906),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_out[22]));
 sky130_fd_sc_hd__buf_2 _11944_ (.A(net907),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_out[23]));
 sky130_fd_sc_hd__buf_2 _11945_ (.A(net908),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_out[24]));
 sky130_fd_sc_hd__buf_2 _11946_ (.A(net909),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_out[25]));
 sky130_fd_sc_hd__buf_2 _11947_ (.A(net910),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_out[26]));
 sky130_fd_sc_hd__buf_2 _11948_ (.A(net911),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_out[27]));
 sky130_fd_sc_hd__buf_2 _11949_ (.A(net912),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_out[28]));
 sky130_fd_sc_hd__buf_2 _11950_ (.A(net913),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_out[29]));
 sky130_fd_sc_hd__buf_2 _11951_ (.A(net914),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_out[30]));
 sky130_fd_sc_hd__buf_2 _11952_ (.A(net915),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_out[31]));
 sky130_fd_sc_hd__buf_2 _11953_ (.A(net916),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_out[32]));
 sky130_fd_sc_hd__buf_2 _11954_ (.A(net917),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_out[33]));
 sky130_fd_sc_hd__conb_1 _10915__918 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(net918));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_0_clk (.A(clknet_4_0_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_Right_102 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_Right_103 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_Right_104 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_Right_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_Right_106 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_Right_107 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_Right_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_Right_109 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_Right_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_Right_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_Right_112 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_Right_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_Right_114 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_Right_115 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_Right_116 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_Right_117 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_Right_118 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_Right_119 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_120 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_121 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_122 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_123 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_124 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_125 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_126 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_127 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_128 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_129 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_130 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_131 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_132 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_134 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_135 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_137 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_140 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_142 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_143 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_144 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_145 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_146 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_147 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_148 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_149 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_150 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_151 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_152 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_153 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_154 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_155 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_156 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_157 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_158 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_159 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_160 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_162 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_163 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_164 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_165 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_166 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_168 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_170 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_171 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_172 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_173 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_174 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_175 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_176 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_177 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_178 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_179 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_180 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_181 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_182 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_183 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_184 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_185 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_186 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_187 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_188 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_190 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_191 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_192 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_194 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_196 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_198 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_199 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_200 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_201 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_202 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_203 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_204 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_205 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_206 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_207 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_208 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_209 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_210 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_211 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_212 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_213 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_214 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_215 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_216 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_217 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_218 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_219 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_220 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_221 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_Left_222 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_Left_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_Left_224 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_Left_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_Left_226 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_Left_227 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_Left_228 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_Left_229 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_Left_230 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_Left_231 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_Left_232 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_Left_233 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_Left_234 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_Left_235 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_Left_236 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_Left_237 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_Left_238 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_Left_239 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_240 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_241 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_242 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_243 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_244 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_245 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_246 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_247 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_248 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_249 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_250 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_251 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_252 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_253 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_254 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_255 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_256 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_257 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_258 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_259 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_260 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_261 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_262 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_263 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_264 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_265 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_266 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_267 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_268 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_269 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_270 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_271 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_272 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_273 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_274 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_275 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_276 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_277 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_278 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_279 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_280 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_281 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_282 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_283 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_284 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_285 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_286 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_287 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_288 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_289 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_290 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_291 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_292 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_293 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_294 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_295 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_296 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_297 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_298 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_299 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_300 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_301 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_302 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_303 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_304 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_305 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_306 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_307 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_308 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_309 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_310 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_311 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_312 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_313 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_314 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_315 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_316 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_317 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_318 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_319 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_320 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_321 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_322 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_323 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_324 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_325 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_326 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_327 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_328 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_329 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_330 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_331 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_332 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_333 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_334 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_335 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_336 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_337 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_338 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_339 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_340 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_341 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_342 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_343 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_344 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_345 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_346 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_347 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_348 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_349 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_350 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_351 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_352 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_353 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_354 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_355 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_356 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_357 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_358 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_359 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_360 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_361 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_362 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_363 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_364 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_365 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_366 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_367 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_368 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_369 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_370 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_371 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_372 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_373 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_374 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_375 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_376 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_377 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_378 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_379 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_380 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_381 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_382 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_383 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_384 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_385 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_386 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_387 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_388 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_389 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_390 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_391 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_392 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_393 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_394 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_395 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_396 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_397 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_398 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_399 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_400 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_401 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_402 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_403 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_404 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_405 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_406 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_407 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_408 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_409 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_410 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_411 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_412 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_413 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_414 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_415 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_416 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_417 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_418 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_419 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_420 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_421 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_422 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_423 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_424 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_425 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_426 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_427 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_428 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_429 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_430 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_431 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_432 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_433 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_434 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_435 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_436 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_437 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_438 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_439 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_440 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_441 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_442 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_443 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_444 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_445 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_446 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_447 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_448 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_449 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_450 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_451 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_452 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_453 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_454 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_455 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_456 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_457 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_458 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_459 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_460 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_461 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_462 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_463 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_464 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_465 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_466 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_467 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_468 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_469 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_470 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_471 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_472 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_473 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_474 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_475 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_476 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_477 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_478 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_479 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_480 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_481 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_482 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_483 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_484 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_485 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_486 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_487 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_488 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_489 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_490 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_491 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_492 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_493 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_494 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_495 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_496 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_497 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_498 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_499 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_500 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_501 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_502 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_503 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_504 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_505 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_506 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_507 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_508 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_509 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_510 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_511 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_512 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_513 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_514 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_515 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_516 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_517 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_518 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_519 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_520 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_521 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_522 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_523 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_524 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_525 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_526 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_527 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_528 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_529 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_530 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_531 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_532 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_533 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_534 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_535 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_536 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_537 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_538 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_539 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_540 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_541 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_542 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_543 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_544 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_545 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_546 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_547 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_548 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_549 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_550 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_551 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_552 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_553 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_554 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_555 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_556 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_557 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_558 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_559 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_560 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_561 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_562 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_563 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_564 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_565 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_566 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_567 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_568 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_569 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_570 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_571 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_572 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_573 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_574 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_575 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_576 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_577 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_578 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_579 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_580 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_581 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_582 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_583 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_584 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_585 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_586 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_587 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_588 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_589 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_590 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_591 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_592 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_593 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_594 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_595 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_596 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_597 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_598 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_599 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_600 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_601 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_602 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_603 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_604 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_605 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_606 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_607 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_608 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_609 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_610 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_611 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_612 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_613 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_614 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_615 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_616 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_617 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_618 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_619 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_620 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_621 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_622 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_623 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_624 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_625 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_626 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_627 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_628 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_629 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_630 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_631 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_632 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_633 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_634 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_635 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_636 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_637 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_638 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_639 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_640 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_641 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_642 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_643 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_644 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_645 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_646 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_647 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_648 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_649 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_650 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_651 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_652 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_653 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_654 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_655 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_656 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_657 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_658 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_659 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_660 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_661 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_662 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_663 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_664 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_665 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_666 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_667 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_668 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_669 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_670 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_671 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_672 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_673 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_674 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_675 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_676 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_677 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_678 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_679 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_680 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_681 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_682 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_683 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_684 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_685 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_686 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_687 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_688 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_689 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_690 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_691 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_692 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_693 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_694 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_695 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_696 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_697 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_698 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_699 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_700 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_701 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_702 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_703 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_704 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_705 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_706 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_707 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_708 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_709 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_710 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_711 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_712 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_713 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_714 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_715 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_716 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_717 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_718 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_719 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_720 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_721 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_722 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_723 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_724 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_725 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_726 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_727 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_728 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_729 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_730 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_731 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_732 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_733 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_734 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_735 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_736 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_737 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_738 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_739 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_740 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_741 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_742 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_743 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_744 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_745 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_746 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_747 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_748 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_749 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_750 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_751 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_752 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_753 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_754 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_755 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_756 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_757 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_758 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_759 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_760 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_761 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_762 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_763 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_764 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_765 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_766 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_767 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_768 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_769 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_770 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_771 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_772 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_773 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_774 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_775 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_776 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_777 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_778 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_779 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_780 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_781 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_782 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_783 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_784 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_785 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_786 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_787 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_788 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_789 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_790 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_791 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_792 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_793 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_794 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_795 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_796 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_797 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_798 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_799 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_800 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_801 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_802 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_803 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_804 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_805 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_806 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_807 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_808 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_809 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_810 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_811 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_812 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_813 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_814 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_815 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_816 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_817 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_818 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_819 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_820 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_821 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_822 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_823 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_824 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_825 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_826 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_827 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_828 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_829 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_830 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_831 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_832 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_833 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_834 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_835 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_836 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_837 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_838 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_839 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_840 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_841 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_842 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_843 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_844 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_845 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_846 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_847 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_848 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_849 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_850 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_851 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_852 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_853 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_854 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_855 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_856 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_857 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_858 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_859 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_860 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_861 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_862 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_863 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_864 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_865 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_866 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_867 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_868 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_869 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_870 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_871 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_872 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_873 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_874 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_875 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_876 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_877 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_878 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_879 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_880 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_881 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_882 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_883 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_884 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_885 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_886 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_887 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_888 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_889 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_890 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_891 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_892 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_893 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_894 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_895 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_896 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_897 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_898 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_899 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_900 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_901 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_902 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_903 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_904 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_905 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_906 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_907 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_908 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_909 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_910 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_911 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_912 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_913 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_914 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_915 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_916 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_917 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_918 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_919 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_920 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_921 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_922 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_923 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_924 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_925 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_926 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_927 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_928 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_929 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_930 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_931 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_932 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_933 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_934 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_935 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_936 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_937 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_938 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_939 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_940 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_941 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_942 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_943 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_944 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_945 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_946 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_947 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_948 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_949 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_950 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_951 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_952 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_953 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_954 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_955 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_956 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_957 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_958 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_959 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_960 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_961 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_962 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_963 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_964 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_965 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_966 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_967 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_968 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_969 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_970 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_971 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_972 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_973 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_974 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_975 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_976 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_977 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_978 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_979 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_980 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_981 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_982 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_983 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_984 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_985 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_986 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_987 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_988 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_989 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_990 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_991 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_992 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_993 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_994 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_995 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_996 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_997 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_998 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_999 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1000 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1001 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1002 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1003 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1004 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1005 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1006 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1007 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1008 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1009 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1010 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1011 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1012 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1013 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1014 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1015 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1016 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1017 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1018 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1019 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1020 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1021 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1022 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1023 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1024 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1025 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1026 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1027 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1028 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1029 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1030 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1031 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1032 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1033 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1034 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1035 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1036 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1037 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1038 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1039 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1040 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1041 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1042 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1043 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1044 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1045 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1046 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1047 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1048 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1049 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1050 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1051 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1052 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1053 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1054 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1055 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1056 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1057 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1058 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1059 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1060 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1061 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1062 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1063 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1064 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1065 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1066 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1067 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1068 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1069 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1070 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1071 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1072 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1073 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1074 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1075 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1076 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1077 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1078 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1079 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1080 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1081 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1082 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1083 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1084 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1085 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1086 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1087 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1088 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1089 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1090 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1091 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1092 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1093 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1094 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1095 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1096 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1097 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1098 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1099 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1100 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1101 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1102 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1103 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1104 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1105 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1106 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1107 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1108 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1109 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1110 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1111 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1112 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1113 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1114 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1115 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1116 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1117 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1118 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1119 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1120 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1121 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1122 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1123 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1124 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1125 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1126 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1127 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1128 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1129 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1130 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1131 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1132 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1133 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1134 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1135 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1136 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1137 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1138 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1139 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1140 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1141 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1142 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1143 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1144 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1145 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1146 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1147 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1148 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1149 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1150 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1151 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1152 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1153 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1154 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1155 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1156 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1157 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1158 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1159 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1160 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1161 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1162 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1163 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1164 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1165 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1166 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1167 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1168 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1169 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1170 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1171 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1172 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1173 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1174 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1175 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1176 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1177 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1178 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1179 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1180 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1181 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1182 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1183 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1184 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1185 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1186 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1187 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1188 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1189 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1190 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1191 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1192 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1193 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1194 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1195 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1196 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1197 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1198 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1199 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1200 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1201 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1202 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1203 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1204 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1205 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1206 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1207 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1208 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1209 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1210 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1211 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1212 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1213 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1214 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1215 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1216 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1217 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1218 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1219 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1220 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1221 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1222 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1223 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1224 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1225 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1226 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1227 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1228 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1229 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1230 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1231 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1232 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1233 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1234 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1235 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1236 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1237 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1238 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1239 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1240 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1241 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1242 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1243 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1244 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1245 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1246 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1247 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1248 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1249 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1250 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1251 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1252 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1253 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1254 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1255 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1256 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1257 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1258 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1259 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1260 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1261 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1262 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1263 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1264 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1265 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1266 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1267 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1268 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1269 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1270 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1271 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1272 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1273 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1274 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1275 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1276 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1277 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1278 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1279 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1280 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1281 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1282 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1283 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1284 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1285 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1286 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1287 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1288 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1289 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1290 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1291 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1292 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1293 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1294 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1295 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1296 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1297 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1298 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1299 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1300 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1301 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1302 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1303 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1304 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1305 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1306 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1307 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1308 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1309 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1310 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1311 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1312 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1313 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1314 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1315 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1316 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1317 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1318 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1319 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1320 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1321 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1322 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1323 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1324 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1325 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1326 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1327 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1328 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1329 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1330 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1331 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1332 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1333 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1334 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1335 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1336 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1337 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1338 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1339 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1340 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1341 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1342 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1343 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1344 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1345 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1346 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1347 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1348 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1349 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1350 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1351 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1352 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1353 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1354 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1355 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1356 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1357 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1358 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1359 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1360 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1361 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1362 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1363 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1364 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1365 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1366 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1367 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1368 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1369 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1370 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1371 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1372 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1373 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1374 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1375 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1376 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1377 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1378 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1379 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1380 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1381 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1382 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1383 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1384 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1385 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1386 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1387 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1388 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1389 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1390 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1391 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1392 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1393 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1394 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1395 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1396 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1397 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1398 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1399 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1400 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1401 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1402 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1403 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1404 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1405 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1406 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1407 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1408 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1409 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1410 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1411 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1412 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1413 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1414 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1415 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1416 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1417 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1418 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1419 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1420 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1421 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1422 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1423 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1424 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1425 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1426 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1427 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1428 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1429 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1430 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1431 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1432 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1433 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1434 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1435 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1436 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1437 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1438 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1439 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1440 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1441 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1442 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1443 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1444 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1445 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1446 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1447 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1448 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1449 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1450 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1451 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1452 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1453 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1454 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1455 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1456 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1457 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1458 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1459 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1460 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1461 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1462 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1463 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1464 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1465 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1466 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1467 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1468 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1469 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1470 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1471 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1472 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1473 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1474 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1475 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1476 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1477 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1478 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1479 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1480 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1481 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1482 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1483 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1484 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1485 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1486 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1487 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1488 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1489 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1490 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1491 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1492 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1493 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1494 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1495 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1496 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1497 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1498 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1499 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1500 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1501 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1502 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1503 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1504 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1505 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1506 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1507 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1508 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1509 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1510 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1511 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1512 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1513 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1514 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1515 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1516 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1517 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1518 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1519 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1520 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1521 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1522 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1523 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1524 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1525 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1526 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1527 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1528 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1529 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1530 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1531 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1532 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1533 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1534 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1535 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1536 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1537 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1538 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1539 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1540 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1541 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1542 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1543 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1544 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1545 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1546 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1547 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1548 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1549 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1550 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1551 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1552 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1553 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1554 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1555 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1556 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1557 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1558 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1559 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1560 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1561 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1562 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1563 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1564 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1565 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1566 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1567 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1568 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1569 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1570 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1571 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1572 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1573 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1574 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1575 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1576 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1577 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1578 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1579 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1580 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1581 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1582 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1583 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1584 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1585 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1586 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1587 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1588 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1589 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1590 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1591 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1592 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1593 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1594 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1595 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1596 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1597 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1598 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1599 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1600 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1601 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1602 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1603 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1604 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1605 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1606 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1607 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1608 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1609 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1610 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1611 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1612 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1613 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1614 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1615 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1616 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1617 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1618 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1619 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1620 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1621 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1622 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1623 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1624 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1625 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1626 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1627 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1628 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1629 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1630 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1631 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1632 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1633 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1634 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1635 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1636 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1637 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1638 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1639 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1640 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1641 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1642 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1643 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1644 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1645 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1646 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1647 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1648 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1649 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1650 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1651 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1652 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1653 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1654 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1655 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1656 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1657 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1658 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1659 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1660 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1661 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1662 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1663 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1664 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1665 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1666 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1667 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1668 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1669 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1670 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1671 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1672 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1673 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1674 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1675 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1676 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1677 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1678 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1679 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1680 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1681 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1682 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1683 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1684 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1685 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1686 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1687 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1688 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1689 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1690 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1691 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1692 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1693 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1694 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1695 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1696 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1697 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1698 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1699 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1700 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1701 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1702 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1703 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1704 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1705 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1706 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1707 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1708 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1709 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1710 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1711 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1712 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1713 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1714 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1715 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1716 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1717 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1718 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1719 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1720 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1721 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1722 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1723 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1724 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1725 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1726 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1727 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1728 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1729 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1730 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1731 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1732 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1733 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1734 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1735 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1736 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1737 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1738 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1739 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1740 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1741 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1742 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1743 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1744 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1745 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1746 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1747 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1748 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1749 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1750 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1751 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1752 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1753 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1754 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1755 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1756 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1757 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1758 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1759 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1760 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1761 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1762 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1763 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1764 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1765 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1766 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1767 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1768 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1769 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1770 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1771 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1772 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1773 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1774 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1775 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1776 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1777 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1778 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1779 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1780 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1781 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1782 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1783 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1784 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1785 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1786 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1787 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1788 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1789 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1790 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1791 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1792 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1793 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1794 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1795 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1796 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1797 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1798 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1799 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1800 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1801 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1802 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1803 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1804 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1805 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1806 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1807 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1808 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1809 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1810 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1811 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1812 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1813 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1814 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1815 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1816 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1817 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1818 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1819 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1820 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1821 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1822 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1823 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1824 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1825 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dlymetal6s2s_1 input1 (.A(ACK_I),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(DAT_I[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(DAT_I[10]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(DAT_I[11]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(DAT_I[12]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(DAT_I[13]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(DAT_I[14]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(DAT_I[15]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(DAT_I[16]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(DAT_I[17]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(DAT_I[18]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(DAT_I[19]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(DAT_I[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(DAT_I[20]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(DAT_I[21]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(DAT_I[22]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(DAT_I[23]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(DAT_I[24]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(DAT_I[25]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(DAT_I[26]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(DAT_I[27]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(DAT_I[28]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(DAT_I[29]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(DAT_I[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(DAT_I[30]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(DAT_I[31]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(DAT_I[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(DAT_I[4]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(DAT_I[5]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(DAT_I[6]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(DAT_I[7]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(DAT_I[8]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(DAT_I[9]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_2 input34 (.A(en),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net34));
 sky130_fd_sc_hd__buf_1 input35 (.A(gpio_in[10]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net35));
 sky130_fd_sc_hd__dlymetal6s2s_1 input36 (.A(gpio_in[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(gpio_in[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net37));
 sky130_fd_sc_hd__buf_1 input38 (.A(gpio_in[4]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net38));
 sky130_fd_sc_hd__buf_1 input39 (.A(gpio_in[5]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net39));
 sky130_fd_sc_hd__buf_1 input40 (.A(gpio_in[6]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net40));
 sky130_fd_sc_hd__buf_1 input41 (.A(gpio_in[7]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net41));
 sky130_fd_sc_hd__buf_1 input42 (.A(gpio_in[8]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net42));
 sky130_fd_sc_hd__buf_1 input43 (.A(gpio_in[9]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_2 input44 (.A(nrst),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net44));
 sky130_fd_sc_hd__buf_2 output45 (.A(net45),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ADR_O[10]));
 sky130_fd_sc_hd__buf_2 output46 (.A(net46),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ADR_O[11]));
 sky130_fd_sc_hd__buf_2 output47 (.A(net47),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ADR_O[12]));
 sky130_fd_sc_hd__buf_2 output48 (.A(net48),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ADR_O[13]));
 sky130_fd_sc_hd__buf_2 output49 (.A(net49),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ADR_O[14]));
 sky130_fd_sc_hd__buf_2 output50 (.A(net50),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ADR_O[15]));
 sky130_fd_sc_hd__buf_2 output51 (.A(net51),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ADR_O[16]));
 sky130_fd_sc_hd__buf_2 output52 (.A(net52),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ADR_O[17]));
 sky130_fd_sc_hd__clkbuf_4 output53 (.A(net53),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ADR_O[18]));
 sky130_fd_sc_hd__buf_2 output54 (.A(net54),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ADR_O[19]));
 sky130_fd_sc_hd__clkbuf_4 output55 (.A(net55),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ADR_O[20]));
 sky130_fd_sc_hd__buf_2 output56 (.A(net56),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ADR_O[21]));
 sky130_fd_sc_hd__buf_2 output57 (.A(net57),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ADR_O[22]));
 sky130_fd_sc_hd__buf_2 output58 (.A(net58),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ADR_O[23]));
 sky130_fd_sc_hd__buf_2 output59 (.A(net59),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ADR_O[24]));
 sky130_fd_sc_hd__buf_2 output60 (.A(net60),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ADR_O[25]));
 sky130_fd_sc_hd__buf_2 output61 (.A(net61),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ADR_O[26]));
 sky130_fd_sc_hd__buf_2 output62 (.A(net62),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ADR_O[28]));
 sky130_fd_sc_hd__buf_2 output63 (.A(net63),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ADR_O[29]));
 sky130_fd_sc_hd__buf_2 output64 (.A(net64),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ADR_O[2]));
 sky130_fd_sc_hd__buf_2 output65 (.A(net65),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ADR_O[3]));
 sky130_fd_sc_hd__buf_2 output66 (.A(net66),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ADR_O[4]));
 sky130_fd_sc_hd__buf_2 output67 (.A(net67),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ADR_O[5]));
 sky130_fd_sc_hd__buf_2 output68 (.A(net68),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ADR_O[6]));
 sky130_fd_sc_hd__buf_2 output69 (.A(net69),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ADR_O[7]));
 sky130_fd_sc_hd__buf_2 output70 (.A(net70),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ADR_O[8]));
 sky130_fd_sc_hd__buf_2 output71 (.A(net71),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ADR_O[9]));
 sky130_fd_sc_hd__buf_2 output72 (.A(net441),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(CYC_O));
 sky130_fd_sc_hd__buf_2 output73 (.A(net73),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(DAT_O[0]));
 sky130_fd_sc_hd__buf_2 output74 (.A(net74),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(DAT_O[10]));
 sky130_fd_sc_hd__buf_2 output75 (.A(net75),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(DAT_O[11]));
 sky130_fd_sc_hd__buf_2 output76 (.A(net76),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(DAT_O[12]));
 sky130_fd_sc_hd__buf_2 output77 (.A(net77),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(DAT_O[13]));
 sky130_fd_sc_hd__buf_2 output78 (.A(net78),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(DAT_O[14]));
 sky130_fd_sc_hd__buf_2 output79 (.A(net79),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(DAT_O[15]));
 sky130_fd_sc_hd__buf_2 output80 (.A(net80),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(DAT_O[16]));
 sky130_fd_sc_hd__buf_2 output81 (.A(net81),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(DAT_O[17]));
 sky130_fd_sc_hd__buf_2 output82 (.A(net82),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(DAT_O[18]));
 sky130_fd_sc_hd__buf_2 output83 (.A(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(DAT_O[19]));
 sky130_fd_sc_hd__buf_2 output84 (.A(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(DAT_O[1]));
 sky130_fd_sc_hd__buf_2 output85 (.A(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(DAT_O[20]));
 sky130_fd_sc_hd__buf_2 output86 (.A(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(DAT_O[21]));
 sky130_fd_sc_hd__buf_2 output87 (.A(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(DAT_O[22]));
 sky130_fd_sc_hd__buf_2 output88 (.A(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(DAT_O[23]));
 sky130_fd_sc_hd__clkbuf_4 output89 (.A(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(DAT_O[24]));
 sky130_fd_sc_hd__buf_2 output90 (.A(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(DAT_O[25]));
 sky130_fd_sc_hd__buf_2 output91 (.A(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(DAT_O[26]));
 sky130_fd_sc_hd__buf_2 output92 (.A(net92),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(DAT_O[27]));
 sky130_fd_sc_hd__clkbuf_4 output93 (.A(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(DAT_O[28]));
 sky130_fd_sc_hd__clkbuf_4 output94 (.A(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(DAT_O[29]));
 sky130_fd_sc_hd__buf_2 output95 (.A(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(DAT_O[2]));
 sky130_fd_sc_hd__clkbuf_4 output96 (.A(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(DAT_O[30]));
 sky130_fd_sc_hd__clkbuf_4 output97 (.A(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(DAT_O[31]));
 sky130_fd_sc_hd__buf_2 output98 (.A(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(DAT_O[3]));
 sky130_fd_sc_hd__buf_2 output99 (.A(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(DAT_O[4]));
 sky130_fd_sc_hd__buf_2 output100 (.A(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(DAT_O[5]));
 sky130_fd_sc_hd__buf_2 output101 (.A(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(DAT_O[6]));
 sky130_fd_sc_hd__buf_2 output102 (.A(net102),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(DAT_O[7]));
 sky130_fd_sc_hd__buf_2 output103 (.A(net103),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(DAT_O[8]));
 sky130_fd_sc_hd__buf_2 output104 (.A(net104),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(DAT_O[9]));
 sky130_fd_sc_hd__buf_2 output105 (.A(net105),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(SEL_O[0]));
 sky130_fd_sc_hd__buf_2 output106 (.A(net106),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(SEL_O[1]));
 sky130_fd_sc_hd__buf_2 output107 (.A(net107),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(SEL_O[2]));
 sky130_fd_sc_hd__buf_2 output108 (.A(net108),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(SEL_O[3]));
 sky130_fd_sc_hd__buf_2 output109 (.A(net109),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(STB_O));
 sky130_fd_sc_hd__buf_2 output110 (.A(net110),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(WE_O));
 sky130_fd_sc_hd__buf_2 output111 (.A(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gpio_out[1]));
 sky130_fd_sc_hd__buf_2 fanout112 (.A(net113),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_4 fanout113 (.A(net114),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_4 fanout114 (.A(_03661_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_4 fanout115 (.A(net116),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_4 fanout116 (.A(_03661_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_4 fanout117 (.A(net122),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_4 fanout118 (.A(net122),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_4 fanout119 (.A(net121),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_4 fanout120 (.A(net121),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net120));
 sky130_fd_sc_hd__buf_2 fanout121 (.A(net122),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_4 fanout122 (.A(_03613_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net122));
 sky130_fd_sc_hd__buf_2 fanout123 (.A(_03612_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net123));
 sky130_fd_sc_hd__buf_1 fanout124 (.A(_03612_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net124));
 sky130_fd_sc_hd__buf_2 fanout125 (.A(net126),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_4 fanout126 (.A(net127),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_4 fanout127 (.A(_03611_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_4 fanout128 (.A(net131),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_4 fanout129 (.A(net130),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_4 fanout130 (.A(net131),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_2 fanout131 (.A(net132),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_2 fanout132 (.A(_03611_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_4 fanout133 (.A(net139),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_2 fanout134 (.A(net139),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net134));
 sky130_fd_sc_hd__buf_2 fanout135 (.A(net138),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_2 fanout136 (.A(net138),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_4 fanout137 (.A(net138),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_4 fanout138 (.A(net139),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net138));
 sky130_fd_sc_hd__buf_2 fanout139 (.A(_03508_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_4 fanout140 (.A(net142),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net140));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout141 (.A(net142),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_2 fanout142 (.A(_03507_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net142));
 sky130_fd_sc_hd__buf_2 fanout143 (.A(net144),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_2 fanout144 (.A(_02909_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_4 fanout145 (.A(net146),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_4 fanout146 (.A(_02909_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_4 fanout147 (.A(_02806_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_4 fanout148 (.A(net149),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_4 fanout149 (.A(net150),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_4 fanout150 (.A(net151),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_4 fanout151 (.A(_03506_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net151));
 sky130_fd_sc_hd__buf_4 fanout152 (.A(net155),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net152));
 sky130_fd_sc_hd__buf_4 fanout153 (.A(net154),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_4 fanout154 (.A(net155),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net154));
 sky130_fd_sc_hd__buf_2 fanout155 (.A(net156),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net155));
 sky130_fd_sc_hd__buf_2 fanout156 (.A(_03506_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net156));
 sky130_fd_sc_hd__buf_4 fanout157 (.A(_03017_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_4 fanout158 (.A(net159),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net158));
 sky130_fd_sc_hd__buf_2 fanout159 (.A(_02908_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net159));
 sky130_fd_sc_hd__buf_2 fanout160 (.A(net161),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net160));
 sky130_fd_sc_hd__buf_2 fanout161 (.A(_02908_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_4 fanout162 (.A(_02805_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_2 fanout163 (.A(_02805_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net163));
 sky130_fd_sc_hd__buf_2 fanout164 (.A(net167),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net164));
 sky130_fd_sc_hd__buf_1 fanout165 (.A(net167),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_4 fanout166 (.A(net167),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net166));
 sky130_fd_sc_hd__buf_2 fanout167 (.A(_02621_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net167));
 sky130_fd_sc_hd__buf_2 fanout168 (.A(net170),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_2 fanout169 (.A(net171),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net169));
 sky130_fd_sc_hd__buf_2 fanout170 (.A(net171),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_4 fanout171 (.A(_02621_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_4 fanout172 (.A(net174),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net172));
 sky130_fd_sc_hd__buf_2 fanout173 (.A(net174),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net173));
 sky130_fd_sc_hd__buf_2 fanout174 (.A(_04616_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net174));
 sky130_fd_sc_hd__buf_2 fanout175 (.A(net177),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net175));
 sky130_fd_sc_hd__buf_2 fanout176 (.A(net177),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_4 fanout177 (.A(_04616_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net177));
 sky130_fd_sc_hd__buf_2 fanout178 (.A(net179),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net178));
 sky130_fd_sc_hd__buf_2 fanout179 (.A(net189),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net179));
 sky130_fd_sc_hd__buf_2 fanout180 (.A(net189),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_2 fanout181 (.A(net189),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net181));
 sky130_fd_sc_hd__buf_2 fanout182 (.A(net185),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net182));
 sky130_fd_sc_hd__buf_2 fanout183 (.A(net185),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net183));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout184 (.A(net185),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net184));
 sky130_fd_sc_hd__buf_1 fanout185 (.A(net189),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net185));
 sky130_fd_sc_hd__buf_2 fanout186 (.A(net188),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net186));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout187 (.A(net188),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net187));
 sky130_fd_sc_hd__buf_2 fanout188 (.A(net189),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net188));
 sky130_fd_sc_hd__clkbuf_2 fanout189 (.A(_04616_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_4 fanout190 (.A(net192),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_2 fanout191 (.A(net192),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net191));
 sky130_fd_sc_hd__buf_2 fanout192 (.A(_04615_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net192));
 sky130_fd_sc_hd__buf_2 fanout193 (.A(net195),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_4 fanout194 (.A(net195),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_4 fanout195 (.A(_04615_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net195));
 sky130_fd_sc_hd__buf_2 fanout196 (.A(net197),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net196));
 sky130_fd_sc_hd__buf_2 fanout197 (.A(net206),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net197));
 sky130_fd_sc_hd__buf_2 fanout198 (.A(net206),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_2 fanout199 (.A(net206),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net199));
 sky130_fd_sc_hd__buf_2 fanout200 (.A(net202),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net200));
 sky130_fd_sc_hd__buf_2 fanout201 (.A(net202),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net201));
 sky130_fd_sc_hd__buf_2 fanout202 (.A(net206),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net202));
 sky130_fd_sc_hd__buf_2 fanout203 (.A(net205),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net203));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout204 (.A(net205),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net204));
 sky130_fd_sc_hd__clkbuf_2 fanout205 (.A(net206),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net205));
 sky130_fd_sc_hd__clkbuf_2 fanout206 (.A(_04615_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net206));
 sky130_fd_sc_hd__clkbuf_4 fanout207 (.A(_02620_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net207));
 sky130_fd_sc_hd__buf_2 fanout208 (.A(_02620_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net208));
 sky130_fd_sc_hd__buf_2 fanout209 (.A(net212),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net209));
 sky130_fd_sc_hd__buf_2 fanout210 (.A(net212),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net210));
 sky130_fd_sc_hd__clkbuf_2 fanout211 (.A(net212),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net211));
 sky130_fd_sc_hd__buf_2 fanout212 (.A(net213),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_4 fanout213 (.A(_02616_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_4 fanout214 (.A(net219),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net214));
 sky130_fd_sc_hd__buf_2 fanout215 (.A(net219),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net215));
 sky130_fd_sc_hd__clkbuf_2 fanout216 (.A(net219),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net216));
 sky130_fd_sc_hd__buf_2 fanout217 (.A(net218),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net217));
 sky130_fd_sc_hd__buf_2 fanout218 (.A(net219),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net218));
 sky130_fd_sc_hd__buf_2 fanout219 (.A(_05254_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net219));
 sky130_fd_sc_hd__buf_2 fanout220 (.A(net223),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net220));
 sky130_fd_sc_hd__clkbuf_4 fanout221 (.A(net223),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net221));
 sky130_fd_sc_hd__clkbuf_2 fanout222 (.A(net223),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net222));
 sky130_fd_sc_hd__clkbuf_2 fanout223 (.A(_05253_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net223));
 sky130_fd_sc_hd__buf_2 fanout224 (.A(net225),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net224));
 sky130_fd_sc_hd__buf_2 fanout225 (.A(net227),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net225));
 sky130_fd_sc_hd__clkbuf_4 fanout226 (.A(net227),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_2 fanout227 (.A(_05253_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net227));
 sky130_fd_sc_hd__clkbuf_4 fanout228 (.A(net229),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net228));
 sky130_fd_sc_hd__clkbuf_4 fanout229 (.A(_05252_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net229));
 sky130_fd_sc_hd__clkbuf_4 fanout230 (.A(net233),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net230));
 sky130_fd_sc_hd__clkbuf_2 fanout231 (.A(net233),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net231));
 sky130_fd_sc_hd__clkbuf_4 fanout232 (.A(net233),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net232));
 sky130_fd_sc_hd__clkbuf_2 fanout233 (.A(_04781_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net233));
 sky130_fd_sc_hd__clkbuf_4 fanout234 (.A(net236),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net234));
 sky130_fd_sc_hd__clkbuf_4 fanout235 (.A(net236),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net235));
 sky130_fd_sc_hd__clkbuf_4 fanout236 (.A(net247),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net236));
 sky130_fd_sc_hd__clkbuf_4 fanout237 (.A(net238),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net237));
 sky130_fd_sc_hd__clkbuf_2 fanout238 (.A(net241),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net238));
 sky130_fd_sc_hd__clkbuf_4 fanout239 (.A(net240),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net239));
 sky130_fd_sc_hd__clkbuf_4 fanout240 (.A(net241),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_2 fanout241 (.A(net247),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net241));
 sky130_fd_sc_hd__clkbuf_4 fanout242 (.A(net243),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net242));
 sky130_fd_sc_hd__clkbuf_4 fanout243 (.A(net246),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net243));
 sky130_fd_sc_hd__clkbuf_4 fanout244 (.A(net246),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net244));
 sky130_fd_sc_hd__buf_2 fanout245 (.A(net246),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net245));
 sky130_fd_sc_hd__buf_2 fanout246 (.A(net247),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net246));
 sky130_fd_sc_hd__clkbuf_2 max_cap247 (.A(_04781_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net247));
 sky130_fd_sc_hd__clkbuf_4 fanout248 (.A(net253),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net248));
 sky130_fd_sc_hd__clkbuf_4 fanout249 (.A(net253),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net249));
 sky130_fd_sc_hd__clkbuf_2 fanout250 (.A(net253),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net250));
 sky130_fd_sc_hd__clkbuf_4 fanout251 (.A(net252),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net251));
 sky130_fd_sc_hd__clkbuf_4 fanout252 (.A(net253),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net252));
 sky130_fd_sc_hd__buf_2 fanout253 (.A(_04337_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net253));
 sky130_fd_sc_hd__buf_2 fanout254 (.A(net255),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net254));
 sky130_fd_sc_hd__clkbuf_2 fanout255 (.A(net256),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net255));
 sky130_fd_sc_hd__clkbuf_2 fanout256 (.A(net259),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net256));
 sky130_fd_sc_hd__buf_2 fanout257 (.A(net259),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net257));
 sky130_fd_sc_hd__clkbuf_2 fanout258 (.A(net259),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net258));
 sky130_fd_sc_hd__clkbuf_2 fanout259 (.A(_04256_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net259));
 sky130_fd_sc_hd__clkbuf_4 fanout260 (.A(_04256_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net260));
 sky130_fd_sc_hd__buf_2 fanout261 (.A(_04256_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net261));
 sky130_fd_sc_hd__buf_2 fanout262 (.A(net263),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net262));
 sky130_fd_sc_hd__buf_2 fanout263 (.A(_04256_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net263));
 sky130_fd_sc_hd__clkbuf_4 fanout264 (.A(net265),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net264));
 sky130_fd_sc_hd__clkbuf_4 fanout265 (.A(_04251_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net265));
 sky130_fd_sc_hd__clkbuf_4 fanout266 (.A(net267),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net266));
 sky130_fd_sc_hd__buf_4 fanout267 (.A(_04251_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net267));
 sky130_fd_sc_hd__clkbuf_4 fanout268 (.A(net270),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net268));
 sky130_fd_sc_hd__clkbuf_2 fanout269 (.A(net270),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net269));
 sky130_fd_sc_hd__clkbuf_4 fanout270 (.A(net273),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net270));
 sky130_fd_sc_hd__clkbuf_4 fanout271 (.A(net272),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net271));
 sky130_fd_sc_hd__clkbuf_4 fanout272 (.A(net273),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net272));
 sky130_fd_sc_hd__clkbuf_2 fanout273 (.A(_03922_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net273));
 sky130_fd_sc_hd__clkbuf_4 fanout274 (.A(net276),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net274));
 sky130_fd_sc_hd__clkbuf_2 fanout275 (.A(net276),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net275));
 sky130_fd_sc_hd__clkbuf_4 fanout276 (.A(net279),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net276));
 sky130_fd_sc_hd__clkbuf_4 fanout277 (.A(net278),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net277));
 sky130_fd_sc_hd__clkbuf_4 fanout278 (.A(net279),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net278));
 sky130_fd_sc_hd__buf_2 fanout279 (.A(_03719_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net279));
 sky130_fd_sc_hd__clkbuf_4 fanout280 (.A(net281),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net280));
 sky130_fd_sc_hd__clkbuf_4 fanout281 (.A(net282),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net281));
 sky130_fd_sc_hd__clkbuf_4 fanout282 (.A(_04249_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net282));
 sky130_fd_sc_hd__buf_4 fanout283 (.A(_04249_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net283));
 sky130_fd_sc_hd__buf_2 fanout284 (.A(_04249_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net284));
 sky130_fd_sc_hd__clkbuf_4 fanout285 (.A(net286),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net285));
 sky130_fd_sc_hd__clkbuf_4 fanout286 (.A(_04249_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net286));
 sky130_fd_sc_hd__buf_2 fanout287 (.A(_03394_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net287));
 sky130_fd_sc_hd__clkbuf_4 fanout288 (.A(_03393_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net288));
 sky130_fd_sc_hd__buf_4 fanout289 (.A(_04111_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net289));
 sky130_fd_sc_hd__buf_2 fanout290 (.A(_04111_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net290));
 sky130_fd_sc_hd__clkbuf_1 max_cap291 (.A(_05185_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net291));
 sky130_fd_sc_hd__clkbuf_4 fanout292 (.A(net295),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net292));
 sky130_fd_sc_hd__clkbuf_4 fanout293 (.A(net294),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net293));
 sky130_fd_sc_hd__clkbuf_4 fanout294 (.A(net295),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net294));
 sky130_fd_sc_hd__buf_2 fanout295 (.A(_04112_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net295));
 sky130_fd_sc_hd__buf_2 fanout296 (.A(_03376_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net296));
 sky130_fd_sc_hd__buf_2 fanout297 (.A(net298),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net297));
 sky130_fd_sc_hd__buf_2 fanout298 (.A(net299),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net298));
 sky130_fd_sc_hd__clkbuf_2 fanout299 (.A(_03244_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net299));
 sky130_fd_sc_hd__buf_4 fanout300 (.A(_03243_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net300));
 sky130_fd_sc_hd__clkbuf_4 fanout301 (.A(_03243_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net301));
 sky130_fd_sc_hd__clkbuf_4 fanout302 (.A(net304),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net302));
 sky130_fd_sc_hd__clkbuf_2 fanout303 (.A(net304),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net303));
 sky130_fd_sc_hd__clkbuf_2 fanout304 (.A(_02918_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net304));
 sky130_fd_sc_hd__clkbuf_4 fanout305 (.A(net306),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net305));
 sky130_fd_sc_hd__buf_2 fanout306 (.A(_02918_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net306));
 sky130_fd_sc_hd__clkbuf_4 fanout307 (.A(net308),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net307));
 sky130_fd_sc_hd__clkbuf_2 fanout308 (.A(_02715_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net308));
 sky130_fd_sc_hd__buf_4 fanout309 (.A(net312),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net309));
 sky130_fd_sc_hd__clkbuf_4 fanout310 (.A(net311),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net310));
 sky130_fd_sc_hd__clkbuf_4 fanout311 (.A(net312),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net311));
 sky130_fd_sc_hd__buf_4 fanout312 (.A(_02606_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net312));
 sky130_fd_sc_hd__clkbuf_4 fanout313 (.A(net317),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net313));
 sky130_fd_sc_hd__clkbuf_2 fanout314 (.A(net317),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net314));
 sky130_fd_sc_hd__clkbuf_4 fanout315 (.A(net317),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net315));
 sky130_fd_sc_hd__clkbuf_2 fanout316 (.A(net317),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net316));
 sky130_fd_sc_hd__clkbuf_2 fanout317 (.A(_05083_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net317));
 sky130_fd_sc_hd__clkbuf_4 fanout318 (.A(net319),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net318));
 sky130_fd_sc_hd__clkbuf_2 fanout319 (.A(net322),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net319));
 sky130_fd_sc_hd__clkbuf_4 fanout320 (.A(net322),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net320));
 sky130_fd_sc_hd__clkbuf_2 fanout321 (.A(net322),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net321));
 sky130_fd_sc_hd__clkbuf_2 fanout322 (.A(_05075_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net322));
 sky130_fd_sc_hd__clkbuf_4 fanout323 (.A(_04917_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net323));
 sky130_fd_sc_hd__clkbuf_4 fanout324 (.A(_04917_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net324));
 sky130_fd_sc_hd__clkbuf_2 fanout325 (.A(_04917_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net325));
 sky130_fd_sc_hd__buf_2 fanout326 (.A(net327),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net326));
 sky130_fd_sc_hd__buf_2 fanout327 (.A(net331),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net327));
 sky130_fd_sc_hd__buf_2 fanout328 (.A(net331),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net328));
 sky130_fd_sc_hd__buf_2 fanout329 (.A(net331),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net329));
 sky130_fd_sc_hd__buf_2 fanout330 (.A(net331),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net330));
 sky130_fd_sc_hd__clkbuf_2 fanout331 (.A(net341),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net331));
 sky130_fd_sc_hd__clkbuf_4 fanout332 (.A(net335),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net332));
 sky130_fd_sc_hd__clkbuf_2 fanout333 (.A(net335),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net333));
 sky130_fd_sc_hd__buf_2 fanout334 (.A(net335),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net334));
 sky130_fd_sc_hd__buf_2 fanout335 (.A(net341),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net335));
 sky130_fd_sc_hd__buf_2 fanout336 (.A(net338),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net336));
 sky130_fd_sc_hd__buf_2 fanout337 (.A(net338),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net337));
 sky130_fd_sc_hd__clkbuf_2 fanout338 (.A(net341),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net338));
 sky130_fd_sc_hd__buf_2 fanout339 (.A(net340),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net339));
 sky130_fd_sc_hd__buf_2 fanout340 (.A(net341),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net340));
 sky130_fd_sc_hd__buf_2 fanout341 (.A(_04637_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net341));
 sky130_fd_sc_hd__clkbuf_4 fanout342 (.A(_04048_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net342));
 sky130_fd_sc_hd__buf_2 fanout343 (.A(_04042_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net343));
 sky130_fd_sc_hd__buf_2 fanout344 (.A(_04042_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net344));
 sky130_fd_sc_hd__clkbuf_4 fanout345 (.A(net346),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net345));
 sky130_fd_sc_hd__buf_2 fanout346 (.A(net348),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net346));
 sky130_fd_sc_hd__clkbuf_4 fanout347 (.A(net348),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net347));
 sky130_fd_sc_hd__buf_2 fanout348 (.A(_02915_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net348));
 sky130_fd_sc_hd__clkbuf_4 fanout349 (.A(net352),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net349));
 sky130_fd_sc_hd__clkbuf_4 fanout350 (.A(net352),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net350));
 sky130_fd_sc_hd__clkbuf_2 fanout351 (.A(net352),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net351));
 sky130_fd_sc_hd__buf_2 fanout352 (.A(net353),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net352));
 sky130_fd_sc_hd__buf_4 fanout353 (.A(_02881_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net353));
 sky130_fd_sc_hd__clkbuf_4 fanout354 (.A(net356),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net354));
 sky130_fd_sc_hd__clkbuf_2 fanout355 (.A(net356),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net355));
 sky130_fd_sc_hd__clkbuf_4 fanout356 (.A(_02609_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net356));
 sky130_fd_sc_hd__buf_2 fanout357 (.A(net358),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net357));
 sky130_fd_sc_hd__clkbuf_4 fanout358 (.A(net359),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net358));
 sky130_fd_sc_hd__buf_4 fanout359 (.A(net360),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net359));
 sky130_fd_sc_hd__buf_4 fanout360 (.A(_02593_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net360));
 sky130_fd_sc_hd__buf_2 fanout361 (.A(_02578_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net361));
 sky130_fd_sc_hd__buf_2 fanout362 (.A(net363),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net362));
 sky130_fd_sc_hd__buf_2 fanout363 (.A(_02571_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net363));
 sky130_fd_sc_hd__buf_2 fanout364 (.A(_02570_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net364));
 sky130_fd_sc_hd__clkbuf_4 fanout365 (.A(net366),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net365));
 sky130_fd_sc_hd__clkbuf_4 fanout366 (.A(_05078_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net366));
 sky130_fd_sc_hd__clkbuf_4 fanout367 (.A(_05077_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net367));
 sky130_fd_sc_hd__buf_2 fanout368 (.A(_05077_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net368));
 sky130_fd_sc_hd__clkbuf_4 fanout369 (.A(net370),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net369));
 sky130_fd_sc_hd__buf_2 fanout370 (.A(_04612_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net370));
 sky130_fd_sc_hd__clkbuf_4 fanout371 (.A(net374),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net371));
 sky130_fd_sc_hd__clkbuf_2 fanout372 (.A(net374),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net372));
 sky130_fd_sc_hd__clkbuf_4 fanout373 (.A(net374),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net373));
 sky130_fd_sc_hd__clkbuf_2 fanout374 (.A(_04612_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net374));
 sky130_fd_sc_hd__buf_2 fanout375 (.A(net376),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net375));
 sky130_fd_sc_hd__buf_2 fanout376 (.A(net386),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net376));
 sky130_fd_sc_hd__buf_2 fanout377 (.A(net386),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net377));
 sky130_fd_sc_hd__clkbuf_2 fanout378 (.A(net386),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net378));
 sky130_fd_sc_hd__buf_2 fanout379 (.A(net382),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net379));
 sky130_fd_sc_hd__buf_2 fanout380 (.A(net382),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net380));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout381 (.A(net382),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net381));
 sky130_fd_sc_hd__buf_1 fanout382 (.A(net386),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net382));
 sky130_fd_sc_hd__buf_2 fanout383 (.A(net385),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net383));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout384 (.A(net385),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net384));
 sky130_fd_sc_hd__buf_2 fanout385 (.A(net386),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net385));
 sky130_fd_sc_hd__clkbuf_2 fanout386 (.A(_04612_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net386));
 sky130_fd_sc_hd__buf_2 fanout387 (.A(net389),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net387));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout388 (.A(net389),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net388));
 sky130_fd_sc_hd__buf_2 fanout389 (.A(net390),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net389));
 sky130_fd_sc_hd__buf_2 fanout390 (.A(net392),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net390));
 sky130_fd_sc_hd__buf_4 fanout391 (.A(net392),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net391));
 sky130_fd_sc_hd__buf_2 fanout392 (.A(_04250_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net392));
 sky130_fd_sc_hd__buf_2 fanout393 (.A(_04049_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net393));
 sky130_fd_sc_hd__buf_4 fanout394 (.A(net397),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net394));
 sky130_fd_sc_hd__buf_4 fanout395 (.A(net396),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net395));
 sky130_fd_sc_hd__buf_4 fanout396 (.A(net397),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net396));
 sky130_fd_sc_hd__clkbuf_4 fanout397 (.A(_02981_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net397));
 sky130_fd_sc_hd__buf_2 fanout398 (.A(net399),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net398));
 sky130_fd_sc_hd__buf_2 fanout399 (.A(net400),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net399));
 sky130_fd_sc_hd__clkbuf_2 fanout400 (.A(net401),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net400));
 sky130_fd_sc_hd__clkbuf_4 fanout401 (.A(_02850_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net401));
 sky130_fd_sc_hd__buf_2 fanout402 (.A(_02810_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net402));
 sky130_fd_sc_hd__clkbuf_2 fanout403 (.A(_02810_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net403));
 sky130_fd_sc_hd__clkbuf_4 fanout404 (.A(_02810_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net404));
 sky130_fd_sc_hd__clkbuf_2 fanout405 (.A(_02810_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net405));
 sky130_fd_sc_hd__clkbuf_4 fanout406 (.A(_02786_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net406));
 sky130_fd_sc_hd__clkbuf_2 fanout407 (.A(_02786_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net407));
 sky130_fd_sc_hd__buf_2 fanout408 (.A(net409),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net408));
 sky130_fd_sc_hd__clkbuf_4 fanout409 (.A(net411),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net409));
 sky130_fd_sc_hd__clkbuf_4 fanout410 (.A(net411),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net410));
 sky130_fd_sc_hd__buf_4 fanout411 (.A(_02611_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net411));
 sky130_fd_sc_hd__clkbuf_2 fanout412 (.A(_02580_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net412));
 sky130_fd_sc_hd__buf_2 fanout413 (.A(net414),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net413));
 sky130_fd_sc_hd__buf_2 fanout414 (.A(_02569_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net414));
 sky130_fd_sc_hd__buf_2 fanout415 (.A(_02568_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net415));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout416 (.A(_02568_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net416));
 sky130_fd_sc_hd__clkbuf_4 fanout417 (.A(net422),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net417));
 sky130_fd_sc_hd__clkbuf_4 fanout418 (.A(net422),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net418));
 sky130_fd_sc_hd__clkbuf_2 fanout419 (.A(net422),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net419));
 sky130_fd_sc_hd__buf_2 fanout420 (.A(net421),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net420));
 sky130_fd_sc_hd__clkbuf_4 fanout421 (.A(net422),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net421));
 sky130_fd_sc_hd__clkbuf_4 fanout422 (.A(_02560_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net422));
 sky130_fd_sc_hd__clkbuf_4 fanout423 (.A(_02555_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net423));
 sky130_fd_sc_hd__clkbuf_2 fanout424 (.A(_02555_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net424));
 sky130_fd_sc_hd__buf_2 fanout425 (.A(net428),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net425));
 sky130_fd_sc_hd__buf_2 fanout426 (.A(net428),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net426));
 sky130_fd_sc_hd__clkbuf_2 fanout427 (.A(net428),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net427));
 sky130_fd_sc_hd__clkbuf_2 fanout428 (.A(_02549_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net428));
 sky130_fd_sc_hd__clkbuf_4 fanout429 (.A(_02548_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net429));
 sky130_fd_sc_hd__buf_2 fanout430 (.A(_02548_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net430));
 sky130_fd_sc_hd__clkbuf_4 fanout431 (.A(net434),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net431));
 sky130_fd_sc_hd__buf_2 fanout432 (.A(net433),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net432));
 sky130_fd_sc_hd__buf_2 fanout433 (.A(net434),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net433));
 sky130_fd_sc_hd__clkbuf_2 fanout434 (.A(_02419_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net434));
 sky130_fd_sc_hd__clkbuf_4 fanout435 (.A(_02419_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net435));
 sky130_fd_sc_hd__buf_2 fanout436 (.A(_02419_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net436));
 sky130_fd_sc_hd__buf_2 fanout437 (.A(net438),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net437));
 sky130_fd_sc_hd__clkbuf_4 fanout438 (.A(_02419_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net438));
 sky130_fd_sc_hd__clkbuf_4 fanout439 (.A(net440),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net439));
 sky130_fd_sc_hd__clkbuf_2 fanout440 (.A(_02404_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net440));
 sky130_fd_sc_hd__clkbuf_4 fanout441 (.A(net72),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net441));
 sky130_fd_sc_hd__buf_2 fanout442 (.A(net443),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net442));
 sky130_fd_sc_hd__buf_2 fanout443 (.A(net444),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net443));
 sky130_fd_sc_hd__clkbuf_4 fanout444 (.A(net72),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net444));
 sky130_fd_sc_hd__buf_2 fanout445 (.A(\top.TRN_char_index[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net445));
 sky130_fd_sc_hd__buf_2 fanout446 (.A(net447),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net446));
 sky130_fd_sc_hd__buf_2 fanout447 (.A(net450),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net447));
 sky130_fd_sc_hd__buf_2 fanout448 (.A(net449),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net448));
 sky130_fd_sc_hd__clkbuf_4 fanout449 (.A(net450),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net449));
 sky130_fd_sc_hd__buf_1 fanout450 (.A(\top.sram_interface.write_HT_fin_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net450));
 sky130_fd_sc_hd__clkbuf_4 fanout451 (.A(net452),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net451));
 sky130_fd_sc_hd__buf_2 fanout452 (.A(\top.controller.state_reg[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net452));
 sky130_fd_sc_hd__clkbuf_4 fanout453 (.A(net454),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net453));
 sky130_fd_sc_hd__clkbuf_4 fanout454 (.A(\top.controller.state_reg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net454));
 sky130_fd_sc_hd__clkbuf_4 fanout455 (.A(net457),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net455));
 sky130_fd_sc_hd__buf_2 fanout456 (.A(net457),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net456));
 sky130_fd_sc_hd__buf_2 fanout457 (.A(\top.controller.state_reg[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net457));
 sky130_fd_sc_hd__buf_2 fanout458 (.A(net459),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net458));
 sky130_fd_sc_hd__clkbuf_4 fanout459 (.A(\top.controller.state_reg[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net459));
 sky130_fd_sc_hd__buf_2 fanout460 (.A(net462),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net460));
 sky130_fd_sc_hd__clkbuf_2 fanout461 (.A(net462),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net461));
 sky130_fd_sc_hd__buf_2 fanout462 (.A(net466),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net462));
 sky130_fd_sc_hd__buf_2 fanout463 (.A(net465),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net463));
 sky130_fd_sc_hd__clkbuf_2 fanout464 (.A(net465),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net464));
 sky130_fd_sc_hd__clkbuf_4 fanout465 (.A(net466),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net465));
 sky130_fd_sc_hd__clkbuf_4 fanout466 (.A(\top.controller.state_reg[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net466));
 sky130_fd_sc_hd__clkbuf_4 fanout467 (.A(net469),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net467));
 sky130_fd_sc_hd__clkbuf_4 fanout468 (.A(net469),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net468));
 sky130_fd_sc_hd__clkbuf_4 fanout469 (.A(\top.controller.state_reg[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net469));
 sky130_fd_sc_hd__buf_2 fanout470 (.A(net471),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net470));
 sky130_fd_sc_hd__clkbuf_2 fanout471 (.A(net480),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net471));
 sky130_fd_sc_hd__clkbuf_2 fanout472 (.A(net474),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net472));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout473 (.A(net474),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net473));
 sky130_fd_sc_hd__buf_2 fanout474 (.A(net475),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net474));
 sky130_fd_sc_hd__buf_2 fanout475 (.A(net480),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net475));
 sky130_fd_sc_hd__buf_2 fanout476 (.A(net480),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net476));
 sky130_fd_sc_hd__clkbuf_2 fanout477 (.A(net480),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net477));
 sky130_fd_sc_hd__clkbuf_2 fanout478 (.A(net480),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net478));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout479 (.A(net480),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net479));
 sky130_fd_sc_hd__clkbuf_4 fanout480 (.A(\top.hTree.state[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net480));
 sky130_fd_sc_hd__buf_2 fanout481 (.A(\top.histogram.init ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net481));
 sky130_fd_sc_hd__buf_2 fanout482 (.A(\top.findLeastValue.histo_index[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net482));
 sky130_fd_sc_hd__clkbuf_4 fanout483 (.A(\top.findLeastValue.histo_index[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net483));
 sky130_fd_sc_hd__buf_2 fanout484 (.A(net485),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net484));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout485 (.A(\top.findLeastValue.histo_index[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net485));
 sky130_fd_sc_hd__buf_2 fanout486 (.A(\top.findLeastValue.histo_index[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net486));
 sky130_fd_sc_hd__buf_2 fanout487 (.A(\top.findLeastValue.histo_index[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net487));
 sky130_fd_sc_hd__buf_2 fanout488 (.A(\top.cb_syn.wait_cycle ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net488));
 sky130_fd_sc_hd__buf_1 fanout489 (.A(\top.cb_syn.wait_cycle ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net489));
 sky130_fd_sc_hd__clkbuf_4 fanout490 (.A(net491),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net490));
 sky130_fd_sc_hd__buf_2 fanout491 (.A(\top.cb_syn.char_found ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net491));
 sky130_fd_sc_hd__clkbuf_4 fanout492 (.A(\top.cb_syn.end_cnt[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net492));
 sky130_fd_sc_hd__buf_2 fanout493 (.A(\top.cb_syn.end_cnt[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net493));
 sky130_fd_sc_hd__clkbuf_4 fanout494 (.A(net495),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net494));
 sky130_fd_sc_hd__clkbuf_4 fanout495 (.A(\top.cb_syn.end_cnt[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net495));
 sky130_fd_sc_hd__clkbuf_4 fanout496 (.A(\top.cb_syn.end_cnt[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net496));
 sky130_fd_sc_hd__buf_2 fanout497 (.A(\top.cb_syn.end_cnt[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net497));
 sky130_fd_sc_hd__clkbuf_4 fanout498 (.A(\top.cb_syn.end_cnt[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net498));
 sky130_fd_sc_hd__clkbuf_4 fanout499 (.A(\top.cb_syn.end_cnt[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net499));
 sky130_fd_sc_hd__buf_4 fanout500 (.A(net501),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net500));
 sky130_fd_sc_hd__buf_4 fanout501 (.A(\top.cb_syn.end_cnt[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net501));
 sky130_fd_sc_hd__clkbuf_4 fanout502 (.A(\top.translation.index[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net502));
 sky130_fd_sc_hd__buf_2 fanout503 (.A(\top.translation.index[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net503));
 sky130_fd_sc_hd__clkbuf_4 fanout504 (.A(net505),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net504));
 sky130_fd_sc_hd__clkbuf_4 fanout505 (.A(\top.translation.index[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net505));
 sky130_fd_sc_hd__clkbuf_4 fanout506 (.A(\top.translation.index[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net506));
 sky130_fd_sc_hd__buf_2 fanout507 (.A(\top.translation.index[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net507));
 sky130_fd_sc_hd__buf_4 fanout508 (.A(net509),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net508));
 sky130_fd_sc_hd__clkbuf_4 fanout509 (.A(net512),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net509));
 sky130_fd_sc_hd__clkbuf_4 fanout510 (.A(net512),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net510));
 sky130_fd_sc_hd__buf_4 fanout511 (.A(net512),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net511));
 sky130_fd_sc_hd__clkbuf_4 fanout512 (.A(\top.translation.index[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net512));
 sky130_fd_sc_hd__buf_2 fanout513 (.A(\top.translation.resEn ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net513));
 sky130_fd_sc_hd__buf_2 fanout514 (.A(\top.cb_syn.curr_state[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net514));
 sky130_fd_sc_hd__buf_2 fanout515 (.A(net516),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net515));
 sky130_fd_sc_hd__buf_2 fanout516 (.A(\top.cb_syn.pulse_first_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net516));
 sky130_fd_sc_hd__buf_2 fanout517 (.A(net518),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net517));
 sky130_fd_sc_hd__clkbuf_2 fanout518 (.A(net520),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net518));
 sky130_fd_sc_hd__clkbuf_4 fanout519 (.A(net520),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net519));
 sky130_fd_sc_hd__clkbuf_2 fanout520 (.A(\top.cb_syn.char_path_n[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net520));
 sky130_fd_sc_hd__buf_2 fanout521 (.A(\top.cb_syn.curr_state[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net521));
 sky130_fd_sc_hd__clkbuf_2 fanout522 (.A(\top.cb_syn.curr_state[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net522));
 sky130_fd_sc_hd__buf_2 fanout523 (.A(\top.cb_syn.curr_state[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net523));
 sky130_fd_sc_hd__buf_2 fanout524 (.A(net525),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net524));
 sky130_fd_sc_hd__buf_2 fanout525 (.A(\top.cb_syn.curr_state[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net525));
 sky130_fd_sc_hd__buf_2 fanout526 (.A(\top.sram_interface.word_cnt[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net526));
 sky130_fd_sc_hd__buf_2 fanout527 (.A(net528),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net527));
 sky130_fd_sc_hd__buf_4 fanout528 (.A(net532),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net528));
 sky130_fd_sc_hd__clkbuf_4 fanout529 (.A(net530),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net529));
 sky130_fd_sc_hd__clkbuf_4 fanout530 (.A(net531),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net530));
 sky130_fd_sc_hd__clkbuf_2 fanout531 (.A(net532),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net531));
 sky130_fd_sc_hd__clkbuf_4 fanout532 (.A(\top.sram_interface.word_cnt[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net532));
 sky130_fd_sc_hd__buf_2 fanout533 (.A(net535),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net533));
 sky130_fd_sc_hd__buf_2 fanout534 (.A(net535),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net534));
 sky130_fd_sc_hd__buf_2 fanout535 (.A(\top.sram_interface.word_cnt[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net535));
 sky130_fd_sc_hd__buf_2 fanout536 (.A(\top.sram_interface.word_cnt[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net536));
 sky130_fd_sc_hd__buf_4 fanout537 (.A(\top.sram_interface.word_cnt[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net537));
 sky130_fd_sc_hd__buf_2 fanout538 (.A(\top.sram_interface.word_cnt[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net538));
 sky130_fd_sc_hd__clkbuf_4 fanout539 (.A(net541),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net539));
 sky130_fd_sc_hd__clkbuf_4 fanout540 (.A(net541),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net540));
 sky130_fd_sc_hd__clkbuf_2 fanout541 (.A(\top.sram_interface.word_cnt[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net541));
 sky130_fd_sc_hd__buf_2 fanout542 (.A(net543),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net542));
 sky130_fd_sc_hd__buf_1 fanout543 (.A(net544),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net543));
 sky130_fd_sc_hd__clkbuf_2 fanout544 (.A(\top.sram_interface.word_cnt[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net544));
 sky130_fd_sc_hd__buf_2 fanout545 (.A(net546),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net545));
 sky130_fd_sc_hd__buf_4 fanout546 (.A(\top.sram_interface.word_cnt[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net546));
 sky130_fd_sc_hd__clkbuf_4 fanout547 (.A(net548),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net547));
 sky130_fd_sc_hd__clkbuf_4 fanout548 (.A(net549),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net548));
 sky130_fd_sc_hd__clkbuf_2 fanout549 (.A(\top.sram_interface.word_cnt[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net549));
 sky130_fd_sc_hd__buf_2 fanout550 (.A(\top.cb_syn.h_element[63] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net550));
 sky130_fd_sc_hd__clkbuf_2 fanout551 (.A(net553),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net551));
 sky130_fd_sc_hd__clkbuf_2 fanout552 (.A(net553),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net552));
 sky130_fd_sc_hd__clkbuf_2 fanout553 (.A(net571),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net553));
 sky130_fd_sc_hd__clkbuf_2 fanout554 (.A(net571),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net554));
 sky130_fd_sc_hd__buf_1 fanout555 (.A(net571),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net555));
 sky130_fd_sc_hd__clkbuf_2 fanout556 (.A(net558),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net556));
 sky130_fd_sc_hd__clkbuf_2 fanout557 (.A(net558),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net557));
 sky130_fd_sc_hd__clkbuf_2 fanout558 (.A(net561),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net558));
 sky130_fd_sc_hd__clkbuf_2 fanout559 (.A(net560),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net559));
 sky130_fd_sc_hd__clkbuf_2 fanout560 (.A(net561),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net560));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout561 (.A(net571),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net561));
 sky130_fd_sc_hd__clkbuf_2 fanout562 (.A(net564),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net562));
 sky130_fd_sc_hd__buf_1 fanout563 (.A(net564),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net563));
 sky130_fd_sc_hd__clkbuf_2 fanout564 (.A(net571),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net564));
 sky130_fd_sc_hd__clkbuf_2 fanout565 (.A(net567),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net565));
 sky130_fd_sc_hd__buf_1 fanout566 (.A(net567),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net566));
 sky130_fd_sc_hd__clkbuf_2 fanout567 (.A(net571),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net567));
 sky130_fd_sc_hd__clkbuf_2 fanout568 (.A(net569),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net568));
 sky130_fd_sc_hd__clkbuf_2 fanout569 (.A(net570),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net569));
 sky130_fd_sc_hd__clkbuf_2 fanout570 (.A(net571),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net570));
 sky130_fd_sc_hd__clkbuf_4 fanout571 (.A(net631),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net571));
 sky130_fd_sc_hd__clkbuf_2 fanout572 (.A(net575),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net572));
 sky130_fd_sc_hd__clkbuf_2 fanout573 (.A(net575),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net573));
 sky130_fd_sc_hd__buf_1 fanout574 (.A(net575),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net574));
 sky130_fd_sc_hd__clkbuf_2 fanout575 (.A(net584),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net575));
 sky130_fd_sc_hd__clkbuf_2 fanout576 (.A(net584),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net576));
 sky130_fd_sc_hd__clkbuf_2 fanout577 (.A(net584),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net577));
 sky130_fd_sc_hd__clkbuf_2 fanout578 (.A(net583),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net578));
 sky130_fd_sc_hd__buf_1 fanout579 (.A(net583),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net579));
 sky130_fd_sc_hd__clkbuf_2 fanout580 (.A(net583),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net580));
 sky130_fd_sc_hd__clkbuf_2 fanout581 (.A(net582),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net581));
 sky130_fd_sc_hd__clkbuf_2 fanout582 (.A(net583),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net582));
 sky130_fd_sc_hd__clkbuf_2 fanout583 (.A(net584),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net583));
 sky130_fd_sc_hd__clkbuf_2 fanout584 (.A(net631),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net584));
 sky130_fd_sc_hd__clkbuf_2 fanout585 (.A(net588),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net585));
 sky130_fd_sc_hd__clkbuf_2 fanout586 (.A(net588),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net586));
 sky130_fd_sc_hd__clkbuf_2 fanout587 (.A(net588),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net587));
 sky130_fd_sc_hd__clkbuf_2 fanout588 (.A(net631),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net588));
 sky130_fd_sc_hd__clkbuf_2 fanout589 (.A(net590),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net589));
 sky130_fd_sc_hd__clkbuf_2 fanout590 (.A(net592),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net590));
 sky130_fd_sc_hd__clkbuf_2 fanout591 (.A(net592),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net591));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout592 (.A(net631),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net592));
 sky130_fd_sc_hd__clkbuf_2 fanout593 (.A(net594),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net593));
 sky130_fd_sc_hd__buf_1 fanout594 (.A(net612),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net594));
 sky130_fd_sc_hd__clkbuf_2 fanout595 (.A(net597),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net595));
 sky130_fd_sc_hd__clkbuf_2 fanout596 (.A(net597),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net596));
 sky130_fd_sc_hd__clkbuf_2 fanout597 (.A(net612),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net597));
 sky130_fd_sc_hd__clkbuf_2 fanout598 (.A(net601),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net598));
 sky130_fd_sc_hd__clkbuf_2 fanout599 (.A(net601),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net599));
 sky130_fd_sc_hd__buf_1 fanout600 (.A(net601),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net600));
 sky130_fd_sc_hd__clkbuf_2 fanout601 (.A(net612),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net601));
 sky130_fd_sc_hd__clkbuf_2 fanout602 (.A(net603),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net602));
 sky130_fd_sc_hd__clkbuf_2 fanout603 (.A(net606),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net603));
 sky130_fd_sc_hd__clkbuf_2 fanout604 (.A(net605),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net604));
 sky130_fd_sc_hd__clkbuf_2 fanout605 (.A(net606),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net605));
 sky130_fd_sc_hd__buf_1 fanout606 (.A(net612),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net606));
 sky130_fd_sc_hd__clkbuf_2 fanout607 (.A(net608),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net607));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout608 (.A(net611),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net608));
 sky130_fd_sc_hd__clkbuf_2 fanout609 (.A(net611),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net609));
 sky130_fd_sc_hd__clkbuf_2 fanout610 (.A(net611),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net610));
 sky130_fd_sc_hd__clkbuf_2 fanout611 (.A(net612),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net611));
 sky130_fd_sc_hd__buf_2 fanout612 (.A(net630),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net612));
 sky130_fd_sc_hd__clkbuf_2 fanout613 (.A(net615),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net613));
 sky130_fd_sc_hd__clkbuf_2 fanout614 (.A(net615),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net614));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout615 (.A(net630),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net615));
 sky130_fd_sc_hd__clkbuf_2 fanout616 (.A(net630),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net616));
 sky130_fd_sc_hd__clkbuf_2 fanout617 (.A(net618),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net617));
 sky130_fd_sc_hd__clkbuf_2 fanout618 (.A(net621),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net618));
 sky130_fd_sc_hd__clkbuf_2 fanout619 (.A(net621),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net619));
 sky130_fd_sc_hd__clkbuf_2 fanout620 (.A(net621),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net620));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout621 (.A(net630),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net621));
 sky130_fd_sc_hd__clkbuf_2 fanout622 (.A(net623),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net622));
 sky130_fd_sc_hd__clkbuf_2 fanout623 (.A(net629),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net623));
 sky130_fd_sc_hd__clkbuf_2 fanout624 (.A(net629),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net624));
 sky130_fd_sc_hd__clkbuf_2 fanout625 (.A(net626),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net625));
 sky130_fd_sc_hd__clkbuf_2 fanout626 (.A(net629),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net626));
 sky130_fd_sc_hd__clkbuf_2 fanout627 (.A(net628),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net627));
 sky130_fd_sc_hd__buf_2 fanout628 (.A(net629),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net628));
 sky130_fd_sc_hd__buf_2 fanout629 (.A(net630),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net629));
 sky130_fd_sc_hd__clkbuf_2 fanout630 (.A(net631),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net630));
 sky130_fd_sc_hd__buf_2 fanout631 (.A(net44),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net631));
 sky130_fd_sc_hd__clkbuf_2 fanout632 (.A(net638),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net632));
 sky130_fd_sc_hd__buf_1 fanout633 (.A(net638),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net633));
 sky130_fd_sc_hd__clkbuf_2 fanout634 (.A(net638),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net634));
 sky130_fd_sc_hd__buf_1 fanout635 (.A(net638),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net635));
 sky130_fd_sc_hd__clkbuf_2 fanout636 (.A(net637),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net636));
 sky130_fd_sc_hd__clkbuf_2 fanout637 (.A(net638),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net637));
 sky130_fd_sc_hd__buf_2 fanout638 (.A(net643),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net638));
 sky130_fd_sc_hd__clkbuf_2 fanout639 (.A(net643),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net639));
 sky130_fd_sc_hd__buf_1 fanout640 (.A(net643),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net640));
 sky130_fd_sc_hd__clkbuf_2 fanout641 (.A(net643),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net641));
 sky130_fd_sc_hd__buf_1 fanout642 (.A(net643),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net642));
 sky130_fd_sc_hd__clkbuf_2 fanout643 (.A(net651),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net643));
 sky130_fd_sc_hd__clkbuf_2 fanout644 (.A(net647),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net644));
 sky130_fd_sc_hd__buf_1 fanout645 (.A(net647),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net645));
 sky130_fd_sc_hd__clkbuf_2 fanout646 (.A(net647),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net646));
 sky130_fd_sc_hd__clkbuf_2 fanout647 (.A(net651),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net647));
 sky130_fd_sc_hd__clkbuf_2 fanout648 (.A(net651),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net648));
 sky130_fd_sc_hd__clkbuf_2 fanout649 (.A(net651),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net649));
 sky130_fd_sc_hd__clkbuf_2 fanout650 (.A(net651),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net650));
 sky130_fd_sc_hd__buf_2 fanout651 (.A(net712),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net651));
 sky130_fd_sc_hd__clkbuf_2 fanout652 (.A(net661),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net652));
 sky130_fd_sc_hd__buf_1 fanout653 (.A(net661),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net653));
 sky130_fd_sc_hd__clkbuf_2 fanout654 (.A(net661),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net654));
 sky130_fd_sc_hd__clkbuf_2 fanout655 (.A(net661),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net655));
 sky130_fd_sc_hd__clkbuf_2 fanout656 (.A(net657),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net656));
 sky130_fd_sc_hd__clkbuf_2 fanout657 (.A(net660),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net657));
 sky130_fd_sc_hd__clkbuf_2 fanout658 (.A(net660),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net658));
 sky130_fd_sc_hd__buf_1 fanout659 (.A(net660),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net659));
 sky130_fd_sc_hd__clkbuf_2 fanout660 (.A(net661),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net660));
 sky130_fd_sc_hd__clkbuf_2 fanout661 (.A(net670),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net661));
 sky130_fd_sc_hd__clkbuf_2 fanout662 (.A(net670),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net662));
 sky130_fd_sc_hd__buf_1 fanout663 (.A(net670),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net663));
 sky130_fd_sc_hd__clkbuf_2 fanout664 (.A(net665),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net664));
 sky130_fd_sc_hd__clkbuf_2 fanout665 (.A(net670),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net665));
 sky130_fd_sc_hd__clkbuf_2 fanout666 (.A(net669),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net666));
 sky130_fd_sc_hd__clkbuf_2 fanout667 (.A(net668),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net667));
 sky130_fd_sc_hd__buf_2 fanout668 (.A(net669),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net668));
 sky130_fd_sc_hd__clkbuf_2 fanout669 (.A(net670),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net669));
 sky130_fd_sc_hd__clkbuf_2 fanout670 (.A(net712),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net670));
 sky130_fd_sc_hd__clkbuf_2 fanout671 (.A(net680),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net671));
 sky130_fd_sc_hd__buf_1 fanout672 (.A(net680),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net672));
 sky130_fd_sc_hd__clkbuf_2 fanout673 (.A(net680),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net673));
 sky130_fd_sc_hd__clkbuf_2 fanout674 (.A(net680),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net674));
 sky130_fd_sc_hd__clkbuf_2 fanout675 (.A(net679),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net675));
 sky130_fd_sc_hd__buf_1 fanout676 (.A(net679),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net676));
 sky130_fd_sc_hd__clkbuf_2 fanout677 (.A(net678),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net677));
 sky130_fd_sc_hd__clkbuf_2 fanout678 (.A(net679),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net678));
 sky130_fd_sc_hd__buf_1 fanout679 (.A(net680),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net679));
 sky130_fd_sc_hd__clkbuf_2 fanout680 (.A(net712),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net680));
 sky130_fd_sc_hd__clkbuf_2 fanout681 (.A(net689),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net681));
 sky130_fd_sc_hd__clkbuf_2 fanout682 (.A(net689),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net682));
 sky130_fd_sc_hd__clkbuf_2 fanout683 (.A(net689),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net683));
 sky130_fd_sc_hd__buf_1 fanout684 (.A(net689),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net684));
 sky130_fd_sc_hd__clkbuf_2 fanout685 (.A(net689),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net685));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout686 (.A(net689),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net686));
 sky130_fd_sc_hd__clkbuf_2 fanout687 (.A(net688),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net687));
 sky130_fd_sc_hd__clkbuf_2 fanout688 (.A(net689),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net688));
 sky130_fd_sc_hd__clkbuf_4 fanout689 (.A(net712),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net689));
 sky130_fd_sc_hd__clkbuf_2 fanout690 (.A(net694),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net690));
 sky130_fd_sc_hd__clkbuf_2 fanout691 (.A(net693),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net691));
 sky130_fd_sc_hd__clkbuf_2 fanout692 (.A(net693),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net692));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout693 (.A(net694),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net693));
 sky130_fd_sc_hd__buf_1 fanout694 (.A(net700),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net694));
 sky130_fd_sc_hd__clkbuf_2 fanout695 (.A(net696),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net695));
 sky130_fd_sc_hd__clkbuf_2 fanout696 (.A(net700),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net696));
 sky130_fd_sc_hd__clkbuf_2 fanout697 (.A(net700),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net697));
 sky130_fd_sc_hd__buf_1 fanout698 (.A(net700),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net698));
 sky130_fd_sc_hd__clkbuf_2 fanout699 (.A(net700),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net699));
 sky130_fd_sc_hd__clkbuf_2 fanout700 (.A(net711),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net700));
 sky130_fd_sc_hd__clkbuf_2 fanout701 (.A(net702),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net701));
 sky130_fd_sc_hd__clkbuf_2 fanout702 (.A(net711),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net702));
 sky130_fd_sc_hd__clkbuf_2 fanout703 (.A(net711),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net703));
 sky130_fd_sc_hd__clkbuf_2 fanout704 (.A(net711),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net704));
 sky130_fd_sc_hd__clkbuf_2 fanout705 (.A(net710),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net705));
 sky130_fd_sc_hd__buf_1 fanout706 (.A(net707),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net706));
 sky130_fd_sc_hd__clkbuf_2 fanout707 (.A(net710),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net707));
 sky130_fd_sc_hd__clkbuf_2 fanout708 (.A(net709),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net708));
 sky130_fd_sc_hd__clkbuf_2 fanout709 (.A(net710),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net709));
 sky130_fd_sc_hd__clkbuf_2 fanout710 (.A(net711),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net710));
 sky130_fd_sc_hd__clkbuf_2 fanout711 (.A(net712),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net711));
 sky130_fd_sc_hd__clkbuf_4 fanout712 (.A(net44),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net712));
 sky130_fd_sc_hd__clkbuf_4 fanout713 (.A(net714),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net713));
 sky130_fd_sc_hd__clkbuf_4 fanout714 (.A(net715),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net714));
 sky130_fd_sc_hd__buf_2 fanout715 (.A(net37),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net715));
 sky130_fd_sc_hd__clkbuf_2 fanout716 (.A(net718),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net716));
 sky130_fd_sc_hd__clkbuf_2 fanout717 (.A(net718),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net717));
 sky130_fd_sc_hd__clkbuf_2 fanout718 (.A(net736),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net718));
 sky130_fd_sc_hd__clkbuf_2 fanout719 (.A(net736),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net719));
 sky130_fd_sc_hd__buf_1 fanout720 (.A(net736),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net720));
 sky130_fd_sc_hd__clkbuf_2 fanout721 (.A(net723),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net721));
 sky130_fd_sc_hd__clkbuf_2 fanout722 (.A(net723),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net722));
 sky130_fd_sc_hd__clkbuf_2 fanout723 (.A(net726),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net723));
 sky130_fd_sc_hd__clkbuf_2 fanout724 (.A(net725),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net724));
 sky130_fd_sc_hd__clkbuf_2 fanout725 (.A(net726),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net725));
 sky130_fd_sc_hd__clkbuf_2 fanout726 (.A(net736),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net726));
 sky130_fd_sc_hd__clkbuf_2 fanout727 (.A(net729),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net727));
 sky130_fd_sc_hd__buf_1 fanout728 (.A(net729),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net728));
 sky130_fd_sc_hd__clkbuf_2 fanout729 (.A(net736),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net729));
 sky130_fd_sc_hd__clkbuf_2 fanout730 (.A(net732),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net730));
 sky130_fd_sc_hd__buf_1 fanout731 (.A(net732),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net731));
 sky130_fd_sc_hd__clkbuf_2 fanout732 (.A(net736),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net732));
 sky130_fd_sc_hd__clkbuf_2 fanout733 (.A(net734),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net733));
 sky130_fd_sc_hd__clkbuf_2 fanout734 (.A(net735),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net734));
 sky130_fd_sc_hd__clkbuf_2 fanout735 (.A(net736),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net735));
 sky130_fd_sc_hd__clkbuf_4 fanout736 (.A(net796),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net736));
 sky130_fd_sc_hd__clkbuf_2 fanout737 (.A(net740),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net737));
 sky130_fd_sc_hd__clkbuf_2 fanout738 (.A(net740),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net738));
 sky130_fd_sc_hd__buf_1 fanout739 (.A(net740),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net739));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout740 (.A(net749),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net740));
 sky130_fd_sc_hd__clkbuf_2 fanout741 (.A(net749),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net741));
 sky130_fd_sc_hd__clkbuf_2 fanout742 (.A(net749),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net742));
 sky130_fd_sc_hd__clkbuf_2 fanout743 (.A(net748),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net743));
 sky130_fd_sc_hd__buf_1 fanout744 (.A(net748),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net744));
 sky130_fd_sc_hd__clkbuf_2 fanout745 (.A(net748),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net745));
 sky130_fd_sc_hd__clkbuf_2 fanout746 (.A(net747),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net746));
 sky130_fd_sc_hd__clkbuf_2 fanout747 (.A(net748),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net747));
 sky130_fd_sc_hd__clkbuf_2 fanout748 (.A(net749),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net748));
 sky130_fd_sc_hd__clkbuf_2 fanout749 (.A(net796),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net749));
 sky130_fd_sc_hd__clkbuf_2 fanout750 (.A(net753),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net750));
 sky130_fd_sc_hd__clkbuf_2 fanout751 (.A(net753),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net751));
 sky130_fd_sc_hd__clkbuf_2 fanout752 (.A(net753),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net752));
 sky130_fd_sc_hd__clkbuf_2 fanout753 (.A(net796),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net753));
 sky130_fd_sc_hd__clkbuf_2 fanout754 (.A(net755),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net754));
 sky130_fd_sc_hd__clkbuf_2 fanout755 (.A(net757),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net755));
 sky130_fd_sc_hd__clkbuf_2 fanout756 (.A(net757),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net756));
 sky130_fd_sc_hd__clkbuf_2 fanout757 (.A(net796),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net757));
 sky130_fd_sc_hd__clkbuf_2 fanout758 (.A(net759),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net758));
 sky130_fd_sc_hd__buf_1 fanout759 (.A(net777),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net759));
 sky130_fd_sc_hd__clkbuf_2 fanout760 (.A(net762),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net760));
 sky130_fd_sc_hd__clkbuf_2 fanout761 (.A(net762),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net761));
 sky130_fd_sc_hd__clkbuf_2 fanout762 (.A(net777),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net762));
 sky130_fd_sc_hd__clkbuf_2 fanout763 (.A(net766),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net763));
 sky130_fd_sc_hd__clkbuf_2 fanout764 (.A(net766),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net764));
 sky130_fd_sc_hd__buf_1 fanout765 (.A(net766),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net765));
 sky130_fd_sc_hd__clkbuf_2 fanout766 (.A(net777),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net766));
 sky130_fd_sc_hd__clkbuf_2 fanout767 (.A(net768),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net767));
 sky130_fd_sc_hd__clkbuf_2 fanout768 (.A(net771),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net768));
 sky130_fd_sc_hd__clkbuf_2 fanout769 (.A(net770),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net769));
 sky130_fd_sc_hd__clkbuf_2 fanout770 (.A(net771),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net770));
 sky130_fd_sc_hd__clkbuf_2 fanout771 (.A(net777),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net771));
 sky130_fd_sc_hd__clkbuf_2 fanout772 (.A(net773),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net772));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout773 (.A(net776),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net773));
 sky130_fd_sc_hd__clkbuf_2 fanout774 (.A(net776),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net774));
 sky130_fd_sc_hd__clkbuf_2 fanout775 (.A(net776),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net775));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout776 (.A(net777),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net776));
 sky130_fd_sc_hd__clkbuf_2 fanout777 (.A(net795),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net777));
 sky130_fd_sc_hd__clkbuf_2 fanout778 (.A(net780),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net778));
 sky130_fd_sc_hd__clkbuf_2 fanout779 (.A(net780),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net779));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout780 (.A(net795),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net780));
 sky130_fd_sc_hd__clkbuf_2 fanout781 (.A(net795),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net781));
 sky130_fd_sc_hd__clkbuf_2 fanout782 (.A(net783),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net782));
 sky130_fd_sc_hd__clkbuf_2 fanout783 (.A(net786),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net783));
 sky130_fd_sc_hd__clkbuf_2 fanout784 (.A(net786),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net784));
 sky130_fd_sc_hd__clkbuf_2 fanout785 (.A(net786),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net785));
 sky130_fd_sc_hd__clkbuf_2 fanout786 (.A(net795),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net786));
 sky130_fd_sc_hd__clkbuf_2 fanout787 (.A(net788),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net787));
 sky130_fd_sc_hd__clkbuf_2 fanout788 (.A(net794),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net788));
 sky130_fd_sc_hd__clkbuf_2 fanout789 (.A(net794),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net789));
 sky130_fd_sc_hd__clkbuf_2 fanout790 (.A(net791),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net790));
 sky130_fd_sc_hd__clkbuf_2 fanout791 (.A(net794),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net791));
 sky130_fd_sc_hd__clkbuf_2 fanout792 (.A(net793),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net792));
 sky130_fd_sc_hd__clkbuf_2 fanout793 (.A(net794),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net793));
 sky130_fd_sc_hd__buf_2 fanout794 (.A(net795),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net794));
 sky130_fd_sc_hd__buf_2 fanout795 (.A(net796),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net795));
 sky130_fd_sc_hd__clkbuf_4 fanout796 (.A(net34),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net796));
 sky130_fd_sc_hd__clkbuf_2 fanout797 (.A(net803),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net797));
 sky130_fd_sc_hd__buf_1 fanout798 (.A(net803),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net798));
 sky130_fd_sc_hd__clkbuf_2 fanout799 (.A(net803),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net799));
 sky130_fd_sc_hd__buf_1 fanout800 (.A(net803),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net800));
 sky130_fd_sc_hd__clkbuf_2 fanout801 (.A(net802),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net801));
 sky130_fd_sc_hd__clkbuf_2 fanout802 (.A(net803),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net802));
 sky130_fd_sc_hd__buf_2 fanout803 (.A(net808),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net803));
 sky130_fd_sc_hd__clkbuf_2 fanout804 (.A(net808),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net804));
 sky130_fd_sc_hd__buf_1 fanout805 (.A(net808),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net805));
 sky130_fd_sc_hd__clkbuf_2 fanout806 (.A(net808),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net806));
 sky130_fd_sc_hd__buf_1 fanout807 (.A(net808),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net807));
 sky130_fd_sc_hd__clkbuf_2 fanout808 (.A(net816),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net808));
 sky130_fd_sc_hd__clkbuf_2 fanout809 (.A(net812),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net809));
 sky130_fd_sc_hd__buf_1 fanout810 (.A(net812),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net810));
 sky130_fd_sc_hd__clkbuf_2 fanout811 (.A(net812),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net811));
 sky130_fd_sc_hd__clkbuf_2 fanout812 (.A(net816),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net812));
 sky130_fd_sc_hd__clkbuf_2 fanout813 (.A(net816),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net813));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout814 (.A(net816),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net814));
 sky130_fd_sc_hd__clkbuf_2 fanout815 (.A(net816),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net815));
 sky130_fd_sc_hd__buf_2 fanout816 (.A(net877),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net816));
 sky130_fd_sc_hd__clkbuf_2 fanout817 (.A(net826),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net817));
 sky130_fd_sc_hd__buf_1 fanout818 (.A(net826),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net818));
 sky130_fd_sc_hd__clkbuf_2 fanout819 (.A(net826),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net819));
 sky130_fd_sc_hd__clkbuf_2 fanout820 (.A(net826),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net820));
 sky130_fd_sc_hd__clkbuf_2 fanout821 (.A(net822),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net821));
 sky130_fd_sc_hd__clkbuf_2 fanout822 (.A(net825),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net822));
 sky130_fd_sc_hd__clkbuf_2 fanout823 (.A(net825),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net823));
 sky130_fd_sc_hd__buf_1 fanout824 (.A(net825),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net824));
 sky130_fd_sc_hd__clkbuf_2 fanout825 (.A(net826),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net825));
 sky130_fd_sc_hd__clkbuf_2 fanout826 (.A(net835),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net826));
 sky130_fd_sc_hd__clkbuf_2 fanout827 (.A(net835),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net827));
 sky130_fd_sc_hd__buf_1 fanout828 (.A(net835),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net828));
 sky130_fd_sc_hd__clkbuf_2 fanout829 (.A(net830),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net829));
 sky130_fd_sc_hd__clkbuf_2 fanout830 (.A(net835),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net830));
 sky130_fd_sc_hd__clkbuf_2 fanout831 (.A(net834),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net831));
 sky130_fd_sc_hd__clkbuf_2 fanout832 (.A(net833),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net832));
 sky130_fd_sc_hd__clkbuf_2 fanout833 (.A(net834),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net833));
 sky130_fd_sc_hd__clkbuf_2 fanout834 (.A(net835),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net834));
 sky130_fd_sc_hd__buf_2 fanout835 (.A(net877),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net835));
 sky130_fd_sc_hd__clkbuf_2 fanout836 (.A(net845),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net836));
 sky130_fd_sc_hd__buf_1 fanout837 (.A(net845),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net837));
 sky130_fd_sc_hd__clkbuf_2 fanout838 (.A(net845),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net838));
 sky130_fd_sc_hd__clkbuf_2 fanout839 (.A(net845),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net839));
 sky130_fd_sc_hd__clkbuf_2 fanout840 (.A(net844),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net840));
 sky130_fd_sc_hd__buf_1 fanout841 (.A(net844),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net841));
 sky130_fd_sc_hd__clkbuf_2 fanout842 (.A(net843),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net842));
 sky130_fd_sc_hd__clkbuf_2 fanout843 (.A(net844),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net843));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout844 (.A(net845),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net844));
 sky130_fd_sc_hd__clkbuf_2 fanout845 (.A(net877),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net845));
 sky130_fd_sc_hd__clkbuf_2 fanout846 (.A(net854),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net846));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout847 (.A(net854),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net847));
 sky130_fd_sc_hd__clkbuf_2 fanout848 (.A(net854),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net848));
 sky130_fd_sc_hd__buf_1 fanout849 (.A(net854),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net849));
 sky130_fd_sc_hd__clkbuf_2 fanout850 (.A(net854),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net850));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout851 (.A(net854),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net851));
 sky130_fd_sc_hd__clkbuf_2 fanout852 (.A(net853),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net852));
 sky130_fd_sc_hd__clkbuf_2 fanout853 (.A(net854),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net853));
 sky130_fd_sc_hd__buf_2 fanout854 (.A(net877),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net854));
 sky130_fd_sc_hd__clkbuf_2 fanout855 (.A(net859),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net855));
 sky130_fd_sc_hd__clkbuf_2 fanout856 (.A(net858),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net856));
 sky130_fd_sc_hd__clkbuf_2 fanout857 (.A(net858),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net857));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout858 (.A(net859),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net858));
 sky130_fd_sc_hd__clkbuf_2 fanout859 (.A(net865),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net859));
 sky130_fd_sc_hd__clkbuf_2 fanout860 (.A(net861),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net860));
 sky130_fd_sc_hd__clkbuf_2 fanout861 (.A(net865),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net861));
 sky130_fd_sc_hd__clkbuf_2 fanout862 (.A(net865),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net862));
 sky130_fd_sc_hd__buf_1 fanout863 (.A(net865),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net863));
 sky130_fd_sc_hd__clkbuf_2 fanout864 (.A(net865),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net864));
 sky130_fd_sc_hd__clkbuf_2 fanout865 (.A(net876),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net865));
 sky130_fd_sc_hd__clkbuf_2 fanout866 (.A(net867),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net866));
 sky130_fd_sc_hd__clkbuf_2 fanout867 (.A(net876),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net867));
 sky130_fd_sc_hd__clkbuf_2 fanout868 (.A(net876),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net868));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout869 (.A(net876),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net869));
 sky130_fd_sc_hd__clkbuf_2 fanout870 (.A(net875),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net870));
 sky130_fd_sc_hd__buf_1 fanout871 (.A(net872),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net871));
 sky130_fd_sc_hd__clkbuf_2 fanout872 (.A(net875),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net872));
 sky130_fd_sc_hd__clkbuf_2 fanout873 (.A(net874),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net873));
 sky130_fd_sc_hd__clkbuf_2 fanout874 (.A(net875),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net874));
 sky130_fd_sc_hd__clkbuf_2 fanout875 (.A(net876),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net875));
 sky130_fd_sc_hd__clkbuf_2 fanout876 (.A(net877),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net876));
 sky130_fd_sc_hd__clkbuf_4 fanout877 (.A(net34),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net877));
 sky130_fd_sc_hd__conb_1 _11875__878 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(net878));
 sky130_fd_sc_hd__conb_1 _11876__879 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(net879));
 sky130_fd_sc_hd__conb_1 _11877__880 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(net880));
 sky130_fd_sc_hd__conb_1 _11878__881 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(net881));
 sky130_fd_sc_hd__conb_1 _11880__882 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(net882));
 sky130_fd_sc_hd__conb_1 _11881__883 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(net883));
 sky130_fd_sc_hd__conb_1 _11888__884 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(net884));
 sky130_fd_sc_hd__conb_1 _11921__885 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(net885));
 sky130_fd_sc_hd__conb_1 _11923__886 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(net886));
 sky130_fd_sc_hd__conb_1 _11924__887 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(net887));
 sky130_fd_sc_hd__conb_1 _11925__888 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(net888));
 sky130_fd_sc_hd__conb_1 _11926__889 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(net889));
 sky130_fd_sc_hd__conb_1 _11927__890 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(net890));
 sky130_fd_sc_hd__conb_1 _11928__891 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(net891));
 sky130_fd_sc_hd__conb_1 _11929__892 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(net892));
 sky130_fd_sc_hd__conb_1 _11930__893 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(net893));
 sky130_fd_sc_hd__conb_1 _11931__894 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(net894));
 sky130_fd_sc_hd__conb_1 _11932__895 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(net895));
 sky130_fd_sc_hd__conb_1 _11933__896 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(net896));
 sky130_fd_sc_hd__conb_1 _11934__897 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(net897));
 sky130_fd_sc_hd__conb_1 _11935__898 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(net898));
 sky130_fd_sc_hd__conb_1 _11936__899 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(net899));
 sky130_fd_sc_hd__conb_1 _11937__900 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(net900));
 sky130_fd_sc_hd__conb_1 _11938__901 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(net901));
 sky130_fd_sc_hd__conb_1 _11939__902 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(net902));
 sky130_fd_sc_hd__conb_1 _11940__903 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(net903));
 sky130_fd_sc_hd__conb_1 _11941__904 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(net904));
 sky130_fd_sc_hd__conb_1 _11942__905 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(net905));
 sky130_fd_sc_hd__conb_1 _11943__906 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(net906));
 sky130_fd_sc_hd__conb_1 _11944__907 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(net907));
 sky130_fd_sc_hd__conb_1 _11945__908 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(net908));
 sky130_fd_sc_hd__conb_1 _11946__909 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(net909));
 sky130_fd_sc_hd__conb_1 _11947__910 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(net910));
 sky130_fd_sc_hd__conb_1 _11948__911 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(net911));
 sky130_fd_sc_hd__conb_1 _11949__912 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(net912));
 sky130_fd_sc_hd__conb_1 _11950__913 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(net913));
 sky130_fd_sc_hd__conb_1 _11951__914 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(net914));
 sky130_fd_sc_hd__conb_1 _11952__915 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(net915));
 sky130_fd_sc_hd__conb_1 _11953__916 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(net916));
 sky130_fd_sc_hd__conb_1 _11954__917 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(net917));
 sky130_fd_sc_hd__conb_1 _11887__919 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(net919));
 sky130_fd_sc_hd__conb_1 _11889__920 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(net920));
 sky130_fd_sc_hd__conb_1 _11890__921 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(net921));
 sky130_fd_sc_hd__conb_1 _11891__922 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(net922));
 sky130_fd_sc_hd__conb_1 _11892__923 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(net923));
 sky130_fd_sc_hd__conb_1 _11893__924 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(net924));
 sky130_fd_sc_hd__conb_1 _11894__925 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(net925));
 sky130_fd_sc_hd__conb_1 _11895__926 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(net926));
 sky130_fd_sc_hd__conb_1 _11896__927 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(net927));
 sky130_fd_sc_hd__conb_1 _11897__928 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(net928));
 sky130_fd_sc_hd__conb_1 _11898__929 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(net929));
 sky130_fd_sc_hd__conb_1 _11899__930 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(net930));
 sky130_fd_sc_hd__conb_1 _11900__931 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(net931));
 sky130_fd_sc_hd__conb_1 _11901__932 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(net932));
 sky130_fd_sc_hd__conb_1 _11902__933 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(net933));
 sky130_fd_sc_hd__conb_1 _11903__934 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(net934));
 sky130_fd_sc_hd__conb_1 _11904__935 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(net935));
 sky130_fd_sc_hd__conb_1 _11905__936 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(net936));
 sky130_fd_sc_hd__conb_1 _11906__937 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(net937));
 sky130_fd_sc_hd__conb_1 _11907__938 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(net938));
 sky130_fd_sc_hd__conb_1 _11908__939 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(net939));
 sky130_fd_sc_hd__conb_1 _11909__940 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(net940));
 sky130_fd_sc_hd__conb_1 _11910__941 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(net941));
 sky130_fd_sc_hd__conb_1 _11911__942 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(net942));
 sky130_fd_sc_hd__conb_1 _11912__943 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(net943));
 sky130_fd_sc_hd__conb_1 _11913__944 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(net944));
 sky130_fd_sc_hd__conb_1 _11914__945 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(net945));
 sky130_fd_sc_hd__conb_1 _11915__946 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(net946));
 sky130_fd_sc_hd__conb_1 _11916__947 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(net947));
 sky130_fd_sc_hd__conb_1 _11917__948 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(net948));
 sky130_fd_sc_hd__conb_1 _11918__949 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(net949));
 sky130_fd_sc_hd__conb_1 _11919__950 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(net950));
 sky130_fd_sc_hd__conb_1 _11920__951 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(net951));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_1_clk (.A(clknet_4_0_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_2_clk (.A(clknet_4_0_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_3_clk (.A(clknet_4_1_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_4_clk (.A(clknet_4_1_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_5_clk (.A(clknet_4_1_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_6_clk (.A(clknet_4_1_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_7_clk (.A(clknet_4_1_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_8_clk (.A(clknet_4_1_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_9_clk (.A(clknet_4_1_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_10_clk (.A(clknet_4_1_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_11_clk (.A(clknet_4_3_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_12_clk (.A(clknet_4_3_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_13_clk (.A(clknet_4_3_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_14_clk (.A(clknet_4_6_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_15_clk (.A(clknet_4_6_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_16_clk (.A(clknet_4_6_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_17_clk (.A(clknet_4_6_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_18_clk (.A(clknet_4_4_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_19_clk (.A(clknet_4_4_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_20_clk (.A(clknet_4_4_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_21_clk (.A(clknet_4_4_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_22_clk (.A(clknet_4_4_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_23_clk (.A(clknet_4_4_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_24_clk (.A(clknet_4_4_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_25_clk (.A(clknet_4_4_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_26_clk (.A(clknet_4_5_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_27_clk (.A(clknet_4_5_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_28_clk (.A(clknet_4_5_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_29_clk (.A(clknet_4_5_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_30_clk (.A(clknet_4_5_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_31_clk (.A(clknet_4_5_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_32_clk (.A(clknet_4_5_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_33_clk (.A(clknet_4_7_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_34_clk (.A(clknet_4_7_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_35_clk (.A(clknet_4_7_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_36_clk (.A(clknet_4_7_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_37_clk (.A(clknet_4_7_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_38_clk (.A(clknet_4_7_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_39_clk (.A(clknet_4_7_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_40_clk (.A(clknet_4_6_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_41_clk (.A(clknet_4_6_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_42_clk (.A(clknet_4_6_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_43_clk (.A(clknet_4_6_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_44_clk (.A(clknet_4_12_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_45_clk (.A(clknet_4_12_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_46_clk (.A(clknet_4_12_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_47_clk (.A(clknet_4_12_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_48_clk (.A(clknet_4_13_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_49_clk (.A(clknet_4_13_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_50_clk (.A(clknet_4_13_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_51_clk (.A(clknet_4_13_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_52_clk (.A(clknet_4_13_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_53_clk (.A(clknet_4_13_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_54_clk (.A(clknet_4_13_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_55_clk (.A(clknet_4_13_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_56_clk (.A(clknet_4_15_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_57_clk (.A(clknet_4_15_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_58_clk (.A(clknet_4_15_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_58_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_59_clk (.A(clknet_4_15_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_59_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_60_clk (.A(clknet_4_15_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_60_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_61_clk (.A(clknet_4_15_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_61_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_62_clk (.A(clknet_4_15_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_62_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_63_clk (.A(clknet_4_14_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_63_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_64_clk (.A(clknet_4_14_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_64_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_65_clk (.A(clknet_4_14_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_65_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_66_clk (.A(clknet_4_14_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_66_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_67_clk (.A(clknet_4_14_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_67_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_68_clk (.A(clknet_4_14_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_68_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_69_clk (.A(clknet_4_14_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_69_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_70_clk (.A(clknet_4_14_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_70_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_71_clk (.A(clknet_4_12_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_71_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_72_clk (.A(clknet_4_12_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_72_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_73_clk (.A(clknet_4_12_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_73_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_74_clk (.A(clknet_4_12_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_74_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_75_clk (.A(clknet_4_9_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_75_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_76_clk (.A(clknet_4_9_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_76_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_77_clk (.A(clknet_4_9_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_77_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_78_clk (.A(clknet_4_9_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_78_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_79_clk (.A(clknet_4_11_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_79_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_80_clk (.A(clknet_4_11_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_80_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_81_clk (.A(clknet_4_11_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_81_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_82_clk (.A(clknet_4_11_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_82_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_83_clk (.A(clknet_4_11_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_83_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_84_clk (.A(clknet_4_11_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_84_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_85_clk (.A(clknet_4_11_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_85_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_86_clk (.A(clknet_4_10_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_86_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_87_clk (.A(clknet_4_10_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_87_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_88_clk (.A(clknet_4_10_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_88_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_89_clk (.A(clknet_4_10_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_89_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_90_clk (.A(clknet_4_10_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_90_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_91_clk (.A(clknet_4_10_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_91_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_92_clk (.A(clknet_4_10_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_92_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_93_clk (.A(clknet_4_10_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_93_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_94_clk (.A(clknet_4_10_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_94_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_95_clk (.A(clknet_4_8_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_95_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_96_clk (.A(clknet_4_8_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_96_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_97_clk (.A(clknet_4_8_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_97_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_98_clk (.A(clknet_4_8_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_98_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_99_clk (.A(clknet_4_8_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_99_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_100_clk (.A(clknet_4_8_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_100_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_101_clk (.A(clknet_4_8_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_101_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_102_clk (.A(clknet_4_9_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_102_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_103_clk (.A(clknet_4_9_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_103_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_104_clk (.A(clknet_4_9_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_104_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_105_clk (.A(clknet_4_3_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_105_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_106_clk (.A(clknet_4_3_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_106_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_107_clk (.A(clknet_4_3_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_107_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_108_clk (.A(clknet_4_2_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_108_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_109_clk (.A(clknet_4_2_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_109_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_110_clk (.A(clknet_4_2_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_110_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_111_clk (.A(clknet_4_2_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_111_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_112_clk (.A(clknet_4_2_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_112_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_113_clk (.A(clknet_4_2_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_113_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_114_clk (.A(clknet_4_2_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_114_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_115_clk (.A(clknet_4_2_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_115_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_116_clk (.A(clknet_4_0_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_116_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_117_clk (.A(clknet_4_0_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_117_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_118_clk (.A(clknet_4_0_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_118_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_119_clk (.A(clknet_4_0_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_119_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_120_clk (.A(clknet_4_0_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_leaf_120_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\top.controller.fin_HG ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\top.HT_fin_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\top.cb_syn.finished ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\top.controller.fin_FLV ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\top.sram_interface.CB_read_counter ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(_02251_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\top.sram_interface.init_counter[22] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\top.sram_interface.init_counter[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\top.hTree.node_reg[53] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\top.sram_interface.init_counter[23] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\top.sram_interface.init_counter[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\top.sram_interface.init_counter[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\top.hTree.node_reg[27] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\top.sram_interface.init_counter[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\top.sram_interface.init_counter[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\top.sram_interface.init_counter[19] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\top.sram_interface.init_counter[21] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\top.hTree.node_reg[45] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\top.sram_interface.init_counter[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\top.sram_interface.init_counter[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\top.sram_interface.init_counter[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\top.hTree.node_reg[32] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\top.hTree.node_reg[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\top.hTree.node_reg[59] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\top.hTree.node_reg[35] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\top.controller.fin_FINISHED ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\top.hTree.node_reg[57] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\top.hTree.node_reg[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\top.hTree.finish_check ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\top.sram_interface.check ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\top.hTree.node_reg[44] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\top.hTree.node_reg[25] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\top.hTree.node_reg[43] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\top.hTree.tree_reg[51] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\top.hTree.node_reg[26] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\top.hTree.node_reg[22] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\top.hTree.node_reg[62] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\top.hTree.node_reg[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\top.hTree.node_reg[58] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(_02310_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\top.hTree.node_reg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\top.hTree.node_reg[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\top.hTree.tree_reg[50] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\top.hTree.node_reg[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\top.hTree.node_reg[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\top.hTree.tree_reg[48] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\top.hTree.node_reg[21] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\top.hTree.node_reg[61] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\top.hTree.closing ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\top.hTree.node_reg[33] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\top.hTree.node_reg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\top.hTree.node_reg[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\top.hTree.state[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(_01786_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\top.hTree.node_reg[23] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(\top.hTree.node_reg[39] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\top.hTree.node_reg[41] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\top.hTree.tree_reg[52] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\top.hTree.tree_reg[49] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\top.hTree.tree_reg[47] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(net55),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(\top.histogram.sram_out[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\top.hTree.node_reg[40] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\top.hTree.node_reg[42] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(\top.hTree.node_reg[34] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(\top.hTree.node_reg[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(net60),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(\top.hTree.node_reg[56] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(\top.hTree.node_reg[36] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(\top.hTree.node_reg[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(\top.hTree.node_reg[52] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(\top.dut.out[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\top.hTree.node_reg[55] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(\top.hTree.node_reg[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(net110),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(\top.hTree.node_reg[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\top.hTree.node_reg[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(\top.hTree.node_reg[60] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\top.hTree.node_reg[51] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(net53),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(net50),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(net56),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\top.histogram.out_of_init ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(\top.hTree.node_reg[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(net57),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(\top.cb_syn.check_right ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\top.hTree.node_reg[50] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\top.hTree.tree_reg[61] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\top.sram_interface.word_cnt[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(_00040_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(net54),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(net51),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(\top.path[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(\top.histogram.sram_out[23] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\top.path[22] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(\top.sram_interface.word_cnt[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(net48),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(\top.hTree.node_reg[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(\top.cb_syn.char_index[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(\top.path[53] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\top.path[37] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(net61),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(\top.path[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(\top.path[23] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(\top.cb_syn.char_path[23] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(\top.path[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(\top.histogram.sram_out[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(\top.path[42] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(\top.path[26] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(\top.cb_syn.char_path[112] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(\top.path[30] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(\top.cb_syn.char_path[110] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(\top.header_synthesis.header[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(\top.path[81] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(\top.hTree.tree_reg[53] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(\top.cb_syn.char_path[46] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(\top.cb_syn.char_path[28] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(\top.path[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(\top.cb_syn.curr_index[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(\top.cb_syn.char_path[53] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(_01536_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(\top.hTree.tree_reg[57] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(\top.cb_syn.char_path[94] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(net69),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(\top.path[39] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(net67),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(\top.path[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(\top.cb_syn.char_path[120] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(\top.cb_syn.char_path[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(\top.header_synthesis.header[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(\top.cb_syn.char_path[92] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(\top.header_synthesis.header[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(\top.path[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1084));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(\top.cb_syn.left ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1085));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(\top.cb_syn.char_path[69] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(\top.cb_syn.char_path[56] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1087));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(\top.cb_syn.char_path[118] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1088));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(\top.cb_syn.char_path[62] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1089));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(\top.cb_syn.char_path[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1090));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(\top.path[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1091));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(\top.hTree.tree_reg[58] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1092));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(net49),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1093));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(\top.cb_syn.char_path[67] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1094));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(\top.path[108] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1095));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(\top.hTree.node_reg[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1096));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(\top.cb_syn.char_path[111] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1097));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(_01594_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1098));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(\top.cb_syn.char_path[119] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1099));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(\top.cb_syn.char_path[63] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(\top.sram_interface.init_counter[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(_02169_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(\top.translation.writeEn ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(\top.cb_syn.char_path[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(\top.histogram.total[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(\top.path[19] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(\top.path[118] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(\top.histogram.sram_out[19] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(\top.hTree.node_reg[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(\top.path[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(\top.cb_syn.char_path[35] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(\top.cb_syn.char_path[80] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(_01563_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(\top.path[27] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(\top.cb_syn.char_path[105] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(\top.path[29] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(\top.path[50] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(\top.histogram.sram_out[28] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(\top.cb_syn.char_path[127] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(\top.cb_syn.char_path[68] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(\top.cb_syn.char_path[51] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(_01534_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(\top.cb_syn.char_path[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(\top.path[83] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(\top.histogram.sram_out[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(\top.histogram.sram_out[25] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(\top.compVal[24] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(\top.cb_syn.char_path[26] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(\top.cb_syn.char_path[50] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(_01533_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(\top.hTree.tree_reg[60] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(\top.cb_syn.char_path[90] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(\top.cb_syn.char_path[115] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(\top.path[111] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(\top.path[126] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(\top.cb_syn.char_path[52] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(_01535_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(\top.path[34] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(\top.cb_syn.char_path[126] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(\top.histogram.sram_out[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(\top.cb_syn.char_path[36] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(\top.path[38] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(\top.findLeastValue.histo_index[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(\top.path[112] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(\top.histogram.sram_out[21] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(\top.path[72] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(\top.header_synthesis.header[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(\top.path[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(\top.cb_syn.char_path[113] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(\top.path[43] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(\top.cb_syn.char_path[55] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(\top.cb_syn.char_path[30] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(\top.cb_syn.char_path[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(\top.path[56] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(\top.histogram.sram_out[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(\top.path[28] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(\top.cb_syn.char_path[47] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(\top.cb_syn.char_path[96] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(\top.path[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(\top.hTree.tree_reg[62] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(\top.cb_syn.char_path[116] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(\top.path[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(\top.cb_syn.char_path[77] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(\top.hTree.nulls[59] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(\top.path[82] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(\top.path[36] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(\top.histogram.sram_out[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(\top.hTree.nulls[53] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(\top.cb_syn.char_path[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(\top.cb_syn.char_path[21] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(\top.path[57] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(\top.header_synthesis.header[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(net64),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(\top.hTree.tree_reg[55] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(\top.cb_syn.char_path[73] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(\top.cb_syn.char_path[70] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(_01553_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(\top.cb_syn.char_path[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(\top.histogram.sram_out[26] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(\top.path[109] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(\top.cb_syn.char_path[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(\top.path[103] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(\top.cb_syn.char_path[83] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(\top.path[59] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(\top.cb_syn.char_path[88] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(\top.path[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(\top.histogram.sram_out[22] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(\top.path[51] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(\top.path[24] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(\top.hTree.tree_reg[56] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(\top.hTree.nulls[58] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(\top.cb_syn.char_path[32] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(\top.path[121] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(\top.hTree.tree_reg[59] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(net81),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(\top.cb_syn.char_path[79] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(\top.cb_syn.char_path[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(_01500_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(\top.path[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(\top.path[40] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(\top.path[115] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(\top.cb_syn.char_path[103] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(net65),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(\top.path[119] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(\top.hTree.nulls[62] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold256 (.A(\top.path[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(\top.path[44] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(\top.cb_syn.char_path[60] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(\top.cb_syn.char_path[108] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(\top.hTree.nulls[54] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(\top.cb_syn.char_path[100] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(_01583_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(\top.path[86] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(\top.cb_syn.char_path[102] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(\top.path[76] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(\top.path[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold268 (.A(\top.path[52] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(\top.cb_syn.char_path[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(\top.cb_syn.char_path[54] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(\top.hTree.nulls[48] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold272 (.A(\top.path[123] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(\top.path[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold274 (.A(\top.cb_syn.char_path[64] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(net59),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold276 (.A(\top.path[55] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(\top.cb_syn.char_path[19] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(\top.hTree.tree_reg[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(\top.cb_syn.char_path[24] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(\top.cb_syn.char_path[84] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(\top.header_synthesis.header[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(net70),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(\top.path[71] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(\top.cb_syn.char_path[86] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(\top.path[47] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold286 (.A(\top.sram_interface.word_cnt[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(\top.cb_syn.char_path[104] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(\top.path[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(\top.path[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold290 (.A(\top.cb_syn.char_path[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold291 (.A(\top.cb_syn.char_path[101] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(\top.path[62] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(\top.hTree.node_reg[54] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold294 (.A(\top.cb_syn.char_path[81] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold295 (.A(_01564_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold296 (.A(\top.header_synthesis.header[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold297 (.A(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold298 (.A(\top.hTree.nulls[60] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold299 (.A(\top.path[67] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(\top.histogram.sram_out[30] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold301 (.A(\top.hTree.node_reg[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold302 (.A(\top.path[77] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold303 (.A(\top.path[87] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold304 (.A(\top.cb_syn.char_path[45] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold305 (.A(\top.path[46] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold306 (.A(\top.path[70] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold307 (.A(\top.path[66] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold308 (.A(\top.path[107] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold309 (.A(\top.hTree.nulls[49] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold310 (.A(net66),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold311 (.A(\top.cb_syn.char_path[87] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold312 (.A(\top.path[113] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold313 (.A(\top.cb_syn.char_path[82] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold314 (.A(\top.path[90] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold315 (.A(\top.cb_syn.char_path[109] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold316 (.A(\top.path[91] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold317 (.A(\top.hTree.nulls[61] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold318 (.A(\top.cb_syn.char_path[85] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold319 (.A(\top.hTree.nulls[46] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold320 (.A(\top.cb_syn.char_path[37] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold321 (.A(\top.cb_syn.char_path[117] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold322 (.A(_01600_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold323 (.A(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold324 (.A(\top.hTree.node_reg[49] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold325 (.A(_02301_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold326 (.A(\top.cb_syn.char_path[114] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold327 (.A(\top.histogram.sram_out[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold328 (.A(\top.path[122] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold329 (.A(\top.cb_syn.char_path[122] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold330 (.A(\top.sram_interface.write_counter_FLV[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold331 (.A(net102),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold332 (.A(\top.path[58] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold333 (.A(\top.cb_syn.char_path[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold334 (.A(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold335 (.A(\top.path[110] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold336 (.A(\top.cb_syn.char_path[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold337 (.A(\top.hTree.node_reg[37] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold338 (.A(\top.path[94] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold339 (.A(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold340 (.A(\top.cb_syn.char_path[58] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold341 (.A(\top.cb_syn.char_path[93] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold342 (.A(_01576_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold343 (.A(\top.path[120] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold344 (.A(\top.cb_syn.char_path[61] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold345 (.A(\top.path[54] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold346 (.A(\top.cb_syn.char_path[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold347 (.A(\top.cb_syn.char_path[38] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold348 (.A(\top.path[48] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold349 (.A(\top.path[114] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold350 (.A(\top.hTree.nulls[63] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold351 (.A(\top.cb_syn.char_path[99] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold352 (.A(\top.cb_syn.char_path[124] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold353 (.A(\top.cb_syn.char_path[22] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold354 (.A(\top.histogram.sram_out[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold355 (.A(\top.path[127] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold356 (.A(net75),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold357 (.A(\top.path[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold358 (.A(\top.cb_syn.char_path[72] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold359 (.A(\top.cb_syn.char_path[48] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold360 (.A(\top.path[106] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold361 (.A(\top.histogram.sram_out[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold362 (.A(\top.hTree.tree_reg[34] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold363 (.A(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold364 (.A(\top.path[102] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold365 (.A(net78),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold366 (.A(\top.cb_syn.char_path[121] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold367 (.A(\top.hTree.tree_reg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold368 (.A(\top.cb_syn.char_path[40] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold369 (.A(\top.cb_syn.char_path[97] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold370 (.A(\top.cb_syn.char_path[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold371 (.A(\top.cb_syn.char_path[44] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold372 (.A(\top.cb_syn.char_path[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold373 (.A(\top.cb_syn.char_path[33] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold374 (.A(\top.dut.out[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold375 (.A(\top.path[21] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold376 (.A(\top.cb_syn.char_path[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold377 (.A(\top.path[125] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold378 (.A(\top.cb_syn.char_path[95] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold379 (.A(_01578_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold380 (.A(\top.hTree.nulls[47] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold381 (.A(\top.path[41] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold382 (.A(\top.cb_syn.char_path[123] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold383 (.A(\top.cb_syn.char_path[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold384 (.A(\top.hTree.nulls[55] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold385 (.A(\top.cb_syn.char_path[57] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold386 (.A(\top.path[25] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold387 (.A(\top.dut.out[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold388 (.A(\top.path[33] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold389 (.A(\top.hTree.nulls[56] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold390 (.A(\top.path[80] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold391 (.A(\top.cb_syn.char_path[25] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold392 (.A(\top.path[32] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold393 (.A(\top.hTree.nulls[57] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold394 (.A(\top.path[75] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold395 (.A(\top.histogram.sram_out[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold396 (.A(\top.cb_syn.char_path[71] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold397 (.A(_01554_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold398 (.A(\top.cb_syn.char_path[39] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold399 (.A(\top.hTree.tree_reg[19] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold400 (.A(_01808_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold401 (.A(\top.path[68] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold402 (.A(\top.histogram.sram_out[24] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold403 (.A(\top.cb_syn.char_path[34] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold404 (.A(_01517_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold405 (.A(\top.hTree.tree_reg[32] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold406 (.A(\top.cb_syn.char_path[41] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold407 (.A(\top.cb_syn.char_path[106] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold408 (.A(net79),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold409 (.A(\top.cb_syn.char_path[42] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold410 (.A(_01525_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold411 (.A(\top.cb_syn.char_path[74] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold412 (.A(\top.hTree.node_reg[19] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold413 (.A(\top.histogram.total[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold414 (.A(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold415 (.A(\top.histogram.sram_out[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold416 (.A(\top.cb_syn.char_path[75] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold417 (.A(\top.cb_syn.char_path[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold418 (.A(\top.path[100] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold419 (.A(\top.cb_syn.char_path[107] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold420 (.A(\top.hTree.tree_reg[63] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold421 (.A(\top.path[124] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold422 (.A(\top.path[98] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold423 (.A(\top.path[89] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold424 (.A(\top.path[60] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold425 (.A(\top.histogram.sram_out[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold426 (.A(\top.path[65] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold427 (.A(\top.WB.curr_state[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold428 (.A(net71),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold429 (.A(\top.path[69] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold430 (.A(\top.path[79] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold431 (.A(\top.path[116] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold432 (.A(net80),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold433 (.A(\top.cb_syn.char_path[27] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold434 (.A(\top.cb_syn.char_path[65] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold435 (.A(_01548_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold436 (.A(\top.cb_syn.char_path[59] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold437 (.A(\top.hist_data_o[23] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold438 (.A(\top.path[88] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold439 (.A(\top.sram_interface.zero_cnt[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold440 (.A(\top.path[49] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold441 (.A(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold442 (.A(\top.path[95] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold443 (.A(\top.path[74] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold444 (.A(\top.hTree.tree_reg[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold445 (.A(_01809_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold446 (.A(net103),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold447 (.A(\top.path[78] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold448 (.A(\top.path[63] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold449 (.A(\top.path[61] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold450 (.A(\top.path[64] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold451 (.A(\top.cb_syn.char_path[43] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold452 (.A(\top.path[117] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold453 (.A(\top.cb_syn.char_path[98] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold454 (.A(\top.hTree.node_reg[48] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold455 (.A(\top.path[101] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold456 (.A(\top.path[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold457 (.A(\top.header_synthesis.header[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold458 (.A(\top.cb_syn.char_path[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold459 (.A(\top.histogram.sram_out[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold460 (.A(net74),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold461 (.A(\top.path[35] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold462 (.A(\top.cb_syn.char_path[125] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold463 (.A(\top.path[93] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold464 (.A(\top.hTree.node_reg[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold465 (.A(\top.cb_syn.char_path[49] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold466 (.A(\top.cb_syn.curr_index[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold467 (.A(\top.path[99] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold468 (.A(\top.path[85] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold469 (.A(\top.cb_syn.char_path[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold470 (.A(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold471 (.A(\top.histogram.total[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold472 (.A(\top.cb_syn.char_path[66] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold473 (.A(_01549_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold474 (.A(\top.hTree.nulls[52] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold475 (.A(\top.cb_syn.char_path[29] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold476 (.A(_01512_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold477 (.A(\top.sram_interface.zero_cnt[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold478 (.A(\top.histogram.sram_out[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold479 (.A(\top.header_synthesis.count[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold480 (.A(\top.hTree.tree_reg[24] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold481 (.A(_01813_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold482 (.A(\top.hTree.tree_reg[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold483 (.A(net63),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold484 (.A(\top.path[84] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold485 (.A(\top.hTree.tree_reg[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold486 (.A(_01804_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold487 (.A(\top.cb_syn.count[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold488 (.A(\top.cb_syn.char_path[91] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold489 (.A(_01574_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold490 (.A(\top.path[45] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold491 (.A(\top.path[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold492 (.A(\top.hTree.tree_reg[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold493 (.A(_01806_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold494 (.A(\top.hTree.nulls[50] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold495 (.A(\top.histogram.state[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold496 (.A(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold497 (.A(\top.histogram.total[29] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold498 (.A(_03345_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold499 (.A(\top.hTree.tree_reg[44] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold500 (.A(_01833_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold501 (.A(net82),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold502 (.A(\top.path[73] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold503 (.A(\top.histogram.sram_out[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold504 (.A(\top.cb_syn.curr_index[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold505 (.A(\top.histogram.total[23] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold506 (.A(\top.hTree.tree_reg[36] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold507 (.A(\top.hTree.tree_reg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold508 (.A(\top.path[104] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold509 (.A(net92),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold510 (.A(\top.histogram.sram_out[29] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold511 (.A(net76),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold512 (.A(\top.cb_syn.count[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold513 (.A(\top.histogram.sram_out[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold514 (.A(_02095_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold515 (.A(net58),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold516 (.A(\top.histogram.sram_out[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold517 (.A(\top.path[92] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold518 (.A(net104),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold519 (.A(\top.cb_syn.cb_length[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold520 (.A(\top.path[97] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold521 (.A(\top.histogram.sram_out[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold522 (.A(net73),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold523 (.A(\top.hTree.tree_reg[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold524 (.A(\top.hTree.node_reg[38] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold525 (.A(\top.FLV_done ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold526 (.A(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold527 (.A(\top.histogram.total[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold528 (.A(\top.histogram.state[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold529 (.A(_00035_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold530 (.A(\top.hist_data_o[25] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold531 (.A(\top.cb_syn.end_cond ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold532 (.A(_01463_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold533 (.A(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold534 (.A(\top.cb_syn.h_element[53] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold535 (.A(\top.hTree.nulls[51] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold536 (.A(\top.histogram.total[26] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold537 (.A(\top.hTree.node_reg[46] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold538 (.A(\top.sram_interface.zero_cnt[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold539 (.A(\top.hTree.tree_reg[30] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold540 (.A(_01819_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold541 (.A(\top.hTree.tree_reg[35] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold542 (.A(\top.hTree.tree_reg[29] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold543 (.A(_01818_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold544 (.A(\top.hTree.tree_reg[28] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold545 (.A(\top.path[105] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold546 (.A(\top.hTree.tree_reg[43] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold547 (.A(\top.histogram.sram_out[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold548 (.A(\top.cb_syn.curr_index[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold549 (.A(\top.cb_syn.curr_index[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold550 (.A(\top.histogram.total[30] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold551 (.A(\top.histogram.total[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold552 (.A(\top.histogram.total[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold553 (.A(_03355_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold554 (.A(\top.histogram.total[28] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold555 (.A(\top.histogram.total[27] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold556 (.A(_03346_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold557 (.A(\top.header_synthesis.count[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold558 (.A(\top.hist_data_o[26] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold559 (.A(\top.hTree.tree_reg[46] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold560 (.A(\top.hTree.state[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold561 (.A(\top.histogram.total[19] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold562 (.A(\top.cb_syn.char_path[78] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold563 (.A(\top.histogram.state[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold564 (.A(\top.cb_syn.state8 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold565 (.A(\top.hTree.node_reg[24] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold566 (.A(\top.histogram.wr_r_en[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold567 (.A(\top.sram_interface.init_counter[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold568 (.A(\top.histogram.total[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold569 (.A(\top.histogram.total[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold570 (.A(_03351_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold571 (.A(\top.hTree.state[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold572 (.A(_00023_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold573 (.A(\top.hist_data_o[28] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold574 (.A(net47),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold575 (.A(\top.hist_data_o[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold576 (.A(\top.histogram.sram_out[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold577 (.A(\top.hist_data_o[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold578 (.A(\top.hist_data_o[29] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold579 (.A(net77),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold580 (.A(\top.histogram.init_edge ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold581 (.A(\top.histogram.total[22] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold582 (.A(\top.path[96] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold583 (.A(\top.hist_data_o[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold584 (.A(\top.hTree.tree_reg[40] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold585 (.A(\top.hist_data_o[22] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold586 (.A(\top.hTree.tree_reg[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold587 (.A(\top.hTree.tree_reg[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold588 (.A(\top.cb_syn.char_path[76] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold589 (.A(_01559_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold590 (.A(\top.cb_syn.left_check ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold591 (.A(\top.hTree.state[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold592 (.A(_00027_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold593 (.A(\top.histogram.total[24] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold594 (.A(_03348_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold595 (.A(\top.hTree.tree_reg[26] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold596 (.A(_01815_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold597 (.A(net46),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold598 (.A(\top.hist_data_o[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold599 (.A(\top.cb_syn.curr_index[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold600 (.A(\top.hTree.tree_reg[23] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold601 (.A(\top.hTree.tree_reg[21] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold602 (.A(_01810_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold603 (.A(\top.cb_syn.char_path[89] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold604 (.A(\top.cb_syn.curr_path[127] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold605 (.A(\top.cb_syn.curr_index[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold606 (.A(\top.hTree.tree_reg[22] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold607 (.A(\top.hTree.tree_reg[27] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold608 (.A(\top.findLeastValue.sum[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold609 (.A(_01802_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold610 (.A(\top.cb_syn.zero_count[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold611 (.A(\top.hist_data_o[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold612 (.A(\top.histogram.total[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold613 (.A(\top.hTree.tree_reg[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold614 (.A(\top.hTree.tree_reg[25] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold615 (.A(_01814_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold616 (.A(\top.hTree.tree_reg[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold617 (.A(_01805_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold618 (.A(\top.hTree.tree_reg[42] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold619 (.A(\top.hTree.tree_reg[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold620 (.A(_01807_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold621 (.A(\top.cb_syn.pulse_first ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold622 (.A(\top.hTree.tree_reg[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold623 (.A(\top.histogram.wr_r_en[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold624 (.A(\top.hist_addr[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold625 (.A(\top.histogram.sram_out[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold626 (.A(\top.hist_data_o[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold627 (.A(\top.histogram.total[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold628 (.A(\top.hTree.tree_reg[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold629 (.A(\top.hTree.node_reg[63] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold630 (.A(\top.sram_interface.word_cnt[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold631 (.A(\top.hTree.tree_reg[45] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold632 (.A(\top.histogram.total[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold633 (.A(\top.hTree.tree_reg[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold634 (.A(\top.hTree.tree_reg[33] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold635 (.A(_01822_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold636 (.A(net52),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold637 (.A(\top.hTree.state[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold638 (.A(\top.hTree.tree_reg[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold639 (.A(_01799_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold640 (.A(\top.histogram.total[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold641 (.A(\top.controller.fin_reg[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold642 (.A(\top.histogram.total[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold643 (.A(\top.hTree.tree_reg[37] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold644 (.A(\top.cb_syn.count[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold645 (.A(\top.histogram.total[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold646 (.A(\top.histogram.total[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold647 (.A(\top.cb_syn.h_element[62] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold648 (.A(\top.hTree.tree_reg[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold649 (.A(\top.hTree.tree_reg[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold650 (.A(_01800_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold651 (.A(\top.histogram.total[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold652 (.A(\top.hTree.tree_reg[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold653 (.A(\top.hTree.state[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold654 (.A(\top.cb_syn.zero_count[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold655 (.A(\top.hist_data_o[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold656 (.A(\top.hTree.tree_reg[38] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold657 (.A(\top.histogram.total[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold658 (.A(_03362_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold659 (.A(\top.hTree.tree_reg[39] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold660 (.A(\top.histogram.total[25] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold661 (.A(\top.hist_addr[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold662 (.A(_01329_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold663 (.A(\top.sram_interface.init_counter[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold664 (.A(\top.findLeastValue.histo_index[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold665 (.A(\top.findLeastValue.sum[23] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold666 (.A(\top.findLeastValue.histo_index[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold667 (.A(\top.hTree.nullSumIndex[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold668 (.A(\top.hTree.tree_reg[54] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold669 (.A(\top.dut.out[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold670 (.A(\top.cb_syn.cb_enable ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold671 (.A(\top.cb_syn.i[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold672 (.A(\top.hist_data_o[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold673 (.A(\top.findLeastValue.sum[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold674 (.A(\top.hist_data_o[21] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold675 (.A(\top.sram_interface.init_counter[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold676 (.A(\top.findLeastValue.sum[24] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold677 (.A(\top.dut.out[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold678 (.A(\top.hTree.node_reg[28] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold679 (.A(\top.findLeastValue.sum[19] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold680 (.A(\top.sram_interface.write_counter_FLV[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold681 (.A(\top.histogram.total[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold682 (.A(\top.sram_interface.write_counter_FLV[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold683 (.A(\top.hist_data_o[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold684 (.A(\top.translation.write_fin ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold685 (.A(\top.compVal[42] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold686 (.A(\top.hTree.state[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold687 (.A(_00020_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold688 (.A(\top.cw1[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold689 (.A(\top.sram_interface.counter_HTREE[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold690 (.A(\top.cb_syn.count[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold691 (.A(\top.cb_syn.zero_count[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold692 (.A(\top.histogram.total[21] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold693 (.A(\top.cw1[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold694 (.A(\top.hTree.tree_reg[41] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold695 (.A(\top.hist_data_o[30] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold696 (.A(\top.cb_syn.end_check ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold697 (.A(\top.findLeastValue.sum[26] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold698 (.A(\top.cb_syn.i[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold699 (.A(\top.compVal[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold700 (.A(\top.compVal[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold701 (.A(\top.header_synthesis.count[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold702 (.A(\top.histogram.sram_out[27] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold703 (.A(\top.compVal[45] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold704 (.A(\top.hTree.nullSumIndex[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold705 (.A(\top.findLeastValue.sum[29] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold706 (.A(\top.hTree.nullSumIndex[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold707 (.A(\top.histogram.state[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold708 (.A(\top.findLeastValue.sum[28] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold709 (.A(\top.cb_syn.num_lefts[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold710 (.A(\top.cb_syn.num_lefts[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold711 (.A(\top.cb_syn.count[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold712 (.A(\top.hist_data_o[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold713 (.A(\top.cw1[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold714 (.A(\top.hTree.node_reg[47] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold715 (.A(\top.cb_syn.zero_count[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold716 (.A(\top.compVal[25] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold717 (.A(\top.histogram.total[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold718 (.A(\top.findLeastValue.sum[25] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold719 (.A(\top.hTree.nullSumIndex[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold720 (.A(\top.cw1[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold721 (.A(\top.hTree.nullSumIndex[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold722 (.A(\top.cb_syn.count[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold723 (.A(\top.header_synthesis.char_added ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold724 (.A(\top.cb_syn.setup ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold725 (.A(\top.findLeastValue.sum[27] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold726 (.A(\top.hTree.state[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold727 (.A(\top.sram_interface.TRN_counter[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold728 (.A(\top.controller.fin_reg[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold729 (.A(\top.findLeastValue.sum[21] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold730 (.A(\top.controller.fin_reg[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold731 (.A(\top.cb_syn.num_lefts[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold732 (.A(\top.findLeastValue.sum[39] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold733 (.A(\top.dut.bits_in_buf[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold734 (.A(\top.hist_addr[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold735 (.A(\top.hist_data_o[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold736 (.A(\top.compVal[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold737 (.A(\top.cb_syn.i[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold738 (.A(\top.hist_data_o[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold739 (.A(\top.sram_interface.counter_HTREE[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold740 (.A(net45),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold741 (.A(\top.cb_syn.char_path_n[53] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold742 (.A(\top.compVal[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold743 (.A(\top.findLeastValue.histo_index[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold744 (.A(\top.hTree.nullSumIndex[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold745 (.A(\top.findLeastValue.sum[37] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold746 (.A(\top.cb_syn.char_path_n[52] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold747 (.A(\top.compVal[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold748 (.A(\top.hTree.wait_cnt ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold749 (.A(\top.compVal[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold750 (.A(\top.compVal[21] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold751 (.A(\top.sram_interface.init_counter[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold752 (.A(\top.cb_syn.zeroes[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold753 (.A(\top.header_synthesis.start ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold754 (.A(\top.findLeastValue.sum[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold755 (.A(\top.findLeastValue.sum[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold756 (.A(\top.findLeastValue.sum[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold757 (.A(\top.cb_syn.zero_count[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold758 (.A(\top.findLeastValue.sum[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold759 (.A(\top.cb_syn.char_path_n[117] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold760 (.A(\top.findLeastValue.wipe_the_char_1 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold761 (.A(\top.compVal[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold762 (.A(\top.cb_syn.zero_count[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold763 (.A(\top.cb_syn.i[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold764 (.A(\top.findLeastValue.sum[33] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold765 (.A(\top.cb_syn.char_path_n[42] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold766 (.A(\top.cb_syn.zeroes[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold767 (.A(\top.hist_data_o[19] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold768 (.A(\top.cb_syn.char_path_n[80] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold769 (.A(\top.cb_syn.char_path_n[83] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold770 (.A(\top.cb_syn.char_path_n[91] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold771 (.A(\top.cb_syn.zeroes[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold772 (.A(\top.cb_syn.cb_length[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold773 (.A(\top.findLeastValue.sum[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold774 (.A(\top.findLeastValue.sum[30] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold775 (.A(\top.cb_syn.zeroes[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold776 (.A(\top.findLeastValue.sum[43] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold777 (.A(\top.hTree.nullSumIndex[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold778 (.A(\top.compVal[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold779 (.A(\top.compVal[43] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold780 (.A(\top.compVal[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold781 (.A(\top.findLeastValue.sum[45] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold782 (.A(\top.findLeastValue.sum[22] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold783 (.A(\top.compVal[28] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold784 (.A(\top.findLeastValue.sum[42] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold785 (.A(\top.cb_syn.char_path_n[81] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold786 (.A(\top.cb_syn.char_path_n[114] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold787 (.A(\top.cb_syn.char_path_n[119] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold788 (.A(\top.header_synthesis.count[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold789 (.A(\top.hist_addr[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold790 (.A(\top.cb_syn.char_path_n[76] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold791 (.A(\top.cw1[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold792 (.A(\top.findLeastValue.sum[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold793 (.A(\top.cb_syn.char_path_n[111] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold794 (.A(\top.cb_syn.char_path_n[63] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold795 (.A(\top.cb_syn.char_path_n[89] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold796 (.A(\top.cb_syn.char_path_n[50] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold797 (.A(\top.sram_interface.init_counter[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold798 (.A(\top.findLeastValue.sum[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold799 (.A(\top.histogram.state[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold800 (.A(\top.cb_syn.char_path_n[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold801 (.A(\top.cb_syn.char_path_n[82] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold802 (.A(\top.compVal[44] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold803 (.A(\top.cb_syn.char_path_n[29] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold804 (.A(\top.cb_syn.char_path_n[113] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold805 (.A(\top.cb_syn.char_path_n[51] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold806 (.A(\top.sram_interface.init_counter[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold807 (.A(\top.hist_addr[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold808 (.A(\top.cb_syn.char_path_n[112] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold809 (.A(\top.hist_data_o[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold810 (.A(\top.sram_interface.counter_HTREE[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold811 (.A(\top.compVal[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold812 (.A(\top.cb_syn.char_path_n[70] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold813 (.A(\top.compVal[39] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold814 (.A(\top.cb_syn.char_path_n[105] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold815 (.A(\top.cb_syn.char_path_n[22] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold816 (.A(\top.cb_syn.char_path_n[84] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold817 (.A(\top.compVal[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold818 (.A(\top.cb_syn.h_element[58] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold819 (.A(\top.cb_syn.char_path_n[100] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold820 (.A(\top.cb_syn.char_path_n[126] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold821 (.A(\top.cb_syn.char_path_n[108] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold822 (.A(\top.cb_syn.char_path_n[69] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold823 (.A(\top.hist_data_o[27] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold824 (.A(\top.compVal[33] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold825 (.A(\top.compVal[23] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold826 (.A(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold827 (.A(\top.controller.fin_reg[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold828 (.A(\top.cw1[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold829 (.A(\top.cb_syn.h_element[56] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold830 (.A(\top.cb_syn.char_path_n[25] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold831 (.A(\top.cb_syn.char_path_n[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold832 (.A(\top.cb_syn.i[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold833 (.A(\top.compVal[22] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold834 (.A(\top.cb_syn.char_path_n[124] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold835 (.A(\top.histogram.state[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold836 (.A(\top.cb_syn.zeroes[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold837 (.A(\top.cb_syn.char_path_n[92] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold838 (.A(\top.findLeastValue.sum[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold839 (.A(\top.hist_data_o[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold840 (.A(\top.findLeastValue.sum[41] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold841 (.A(\top.cb_syn.char_path_n[75] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold842 (.A(\top.compVal[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold843 (.A(\top.cb_syn.char_path_n[94] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold844 (.A(\top.hTree.node_reg[29] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold845 (.A(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold846 (.A(\top.hist_addr[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold847 (.A(\top.histogram.total[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold848 (.A(\top.hTree.node_reg[60] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold849 (.A(\top.findLeastValue.sum[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold850 (.A(\top.findLeastValue.sum[28] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold851 (.A(\top.compVal[45] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold852 (.A(\top.histogram.total[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold853 (.A(\top.compVal[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold854 (.A(\top.cb_syn.char_path_n[94] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold855 (.A(\top.findLeastValue.sum[23] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold856 (.A(\top.findLeastValue.sum[22] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold857 (.A(\top.cb_syn.char_path_n[89] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1808));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(ACK_I),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(DAT_I[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(DAT_I[10]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(DAT_I[11]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(DAT_I[12]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(DAT_I[13]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(DAT_I[14]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(DAT_I[15]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(DAT_I[16]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(DAT_I[17]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(DAT_I[18]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(DAT_I[19]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(DAT_I[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(DAT_I[20]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(DAT_I[21]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(DAT_I[22]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(DAT_I[23]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(DAT_I[24]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(DAT_I[25]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(DAT_I[26]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(DAT_I[27]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(DAT_I[28]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(DAT_I[29]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(DAT_I[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(DAT_I[30]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(DAT_I[31]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(DAT_I[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(DAT_I[4]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(DAT_I[5]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(DAT_I[6]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(DAT_I[7]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(DAT_I[8]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(DAT_I[9]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout438_A (.DIODE(_02419_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout436_A (.DIODE(_02419_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout435_A (.DIODE(_02419_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout434_A (.DIODE(_02419_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08655__A1 (.DIODE(_02538_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08649__A1 (.DIODE(_02538_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08568__A0 (.DIODE(_02538_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08566__A1 (.DIODE(_02538_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08150__A (.DIODE(_02538_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05903__B (.DIODE(_02538_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08656__A (.DIODE(_02540_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08638__C1 (.DIODE(_02540_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08623__A1 (.DIODE(_02540_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08597__C1 (.DIODE(_02540_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08588__C1 (.DIODE(_02540_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08634__C1 (.DIODE(_02541_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08630__S (.DIODE(_02541_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08618__A (.DIODE(_02541_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08609__B1 (.DIODE(_02541_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08605__A1 (.DIODE(_02541_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08593__B1 (.DIODE(_02541_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08584__B1 (.DIODE(_02541_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08579__B1 (.DIODE(_02541_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08634__A1 (.DIODE(_02542_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08626__S (.DIODE(_02542_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08617__S (.DIODE(_02542_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08610__A1 (.DIODE(_02542_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08602__A (.DIODE(_02542_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08600__S (.DIODE(_02542_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08591__A (.DIODE(_02542_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08582__A (.DIODE(_02542_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08577__A (.DIODE(_02542_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08827__A1 (.DIODE(_02547_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08802__C1 (.DIODE(_02547_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08798__C1 (.DIODE(_02547_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08793__A1 (.DIODE(_02547_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08779__A1 (.DIODE(_02547_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08776__C1 (.DIODE(_02547_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08770__A (.DIODE(_02547_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08768__A (.DIODE(_02547_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08756__C1 (.DIODE(_02547_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09072__B (.DIODE(_02562_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08017__A1 (.DIODE(_02562_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07026__B1 (.DIODE(_02562_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06965__A (.DIODE(_02562_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06597__A2 (.DIODE(_02562_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06596__A (.DIODE(_02562_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05865__A2 (.DIODE(_02562_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05862__B (.DIODE(_02562_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05759__C1 (.DIODE(_02562_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05751__B (.DIODE(_02562_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05762__A (.DIODE(_02564_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05761__B1 (.DIODE(_02564_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09099__A3 (.DIODE(_02582_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05521__B (.DIODE(_02582_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05498__A2 (.DIODE(_02582_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09155__C1 (.DIODE(_02607_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06352__A2 (.DIODE(_02607_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06329__B1 (.DIODE(_02607_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06291__B2 (.DIODE(_02607_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06258__C (.DIODE(_02607_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06241__A1 (.DIODE(_02607_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06195__B2 (.DIODE(_02607_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06166__A3 (.DIODE(_02607_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05523__C1 (.DIODE(_02607_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout208_A (.DIODE(_02620_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout207_A (.DIODE(_02620_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout171_A (.DIODE(_02621_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout167_A (.DIODE(_02621_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05567__B1 (.DIODE(_02644_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05568__B1 (.DIODE(_02646_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05574__B1 (.DIODE(_02651_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05579__B1 (.DIODE(_02654_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05580__B1 (.DIODE(_02656_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05591__B1 (.DIODE(_02664_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05592__B1 (.DIODE(_02666_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05597__B1 (.DIODE(_02669_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05598__B1 (.DIODE(_02671_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05651__A2 (.DIODE(_02714_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout308_A (.DIODE(_02715_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09071__A (.DIODE(_02715_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05657__B1 (.DIODE(_02720_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05663__B1 (.DIODE(_02725_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05670__B1 (.DIODE(_02730_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05675__B1 (.DIODE(_02735_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05705__B1 (.DIODE(_02760_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05711__B1 (.DIODE(_02765_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05717__B1 (.DIODE(_02770_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05724__B1 (.DIODE(_02775_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05729__B1 (.DIODE(_02780_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout163_A (.DIODE(_02805_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout162_A (.DIODE(_02805_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout147_A (.DIODE(_02806_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05765__B1 (.DIODE(_02806_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05764__B1 (.DIODE(_02806_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05768__B1 (.DIODE(_02806_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05767__B1 (.DIODE(_02806_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout405_A (.DIODE(_02810_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout404_A (.DIODE(_02810_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout403_A (.DIODE(_02810_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout402_A (.DIODE(_02810_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05963__C (.DIODE(_02898_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05919__B (.DIODE(_02898_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05918__B (.DIODE(_02898_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09132__A_N (.DIODE(_02906_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05929__A (.DIODE(_02906_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05927__S (.DIODE(_02906_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout161_A (.DIODE(_02908_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout159_A (.DIODE(_02908_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout348_A (.DIODE(_02915_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09071__C_N (.DIODE(_02915_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout306_A (.DIODE(_02918_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout304_A (.DIODE(_02918_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout157_A (.DIODE(_03017_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06139__B1 (.DIODE(_03017_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06140__B1 (.DIODE(_03017_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout301_A (.DIODE(_03243_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout300_A (.DIODE(_03243_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06442__S (.DIODE(_03243_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06434__S (.DIODE(_03243_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout299_A (.DIODE(_03244_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09121__B1 (.DIODE(_03244_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout287_A (.DIODE(_03394_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06910__A (.DIODE(_03394_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06815__A (.DIODE(_03394_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07043__A (.DIODE(_03394_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06614__D (.DIODE(_03411_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06958__B (.DIODE(_03609_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06812__B (.DIODE(_03609_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout132_A (.DIODE(_03611_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout127_A (.DIODE(_03611_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07401__A2 (.DIODE(_03611_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07428__B1 (.DIODE(_03660_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07427__B1 (.DIODE(_03660_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07426__B1 (.DIODE(_03660_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07425__B1 (.DIODE(_03660_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07424__B1 (.DIODE(_03660_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07423__B1 (.DIODE(_03660_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07422__B1 (.DIODE(_03660_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06987__B1 (.DIODE(_03660_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout116_A (.DIODE(_03661_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout114_A (.DIODE(_03661_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07403__A (.DIODE(_03662_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07400__B1 (.DIODE(_03662_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07000__B1 (.DIODE(_03662_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06998__B1 (.DIODE(_03662_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06996__B1 (.DIODE(_03662_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06994__B1 (.DIODE(_03662_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06992__B1 (.DIODE(_03662_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06990__B1 (.DIODE(_03662_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06988__B1 (.DIODE(_03662_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06959__B1 (.DIODE(_03662_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07026__A1 (.DIODE(_03691_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07246__B (.DIODE(_03718_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07043__B (.DIODE(_03718_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07351__A (.DIODE(_03855_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07323__A1 (.DIODE(_03855_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07197__A1 (.DIODE(_03855_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07188__A1 (.DIODE(_03855_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07351__B (.DIODE(_03858_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07323__A2 (.DIODE(_03858_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07197__A2 (.DIODE(_03858_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07188__A2 (.DIODE(_03858_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07256__B2 (.DIODE(_03928_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07262__B2 (.DIODE(_03932_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07572__S (.DIODE(_04110_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07565__S (.DIODE(_04110_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07557__S (.DIODE(_04110_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07550__S (.DIODE(_04110_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07541__S (.DIODE(_04110_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07534__S (.DIODE(_04110_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07526__S (.DIODE(_04110_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07519__S (.DIODE(_04110_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout290_A (.DIODE(_04111_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout289_A (.DIODE(_04111_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07527__A0 (.DIODE(_04119_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07542__A0 (.DIODE(_04134_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07573__A0 (.DIODE(_04165_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07593__B (.DIODE(_04175_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07576__B (.DIODE(_04175_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07653__S (.DIODE(_04212_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07648__S (.DIODE(_04212_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07641__S (.DIODE(_04212_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07634__S (.DIODE(_04212_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07627__S (.DIODE(_04212_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07621__S (.DIODE(_04212_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07614__S (.DIODE(_04212_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07715__S (.DIODE(_04248_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07706__B (.DIODE(_04248_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07700__B (.DIODE(_04248_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07694__B (.DIODE(_04248_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07688__B (.DIODE(_04248_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07682__B (.DIODE(_04248_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07676__B (.DIODE(_04248_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07672__S (.DIODE(_04248_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07668__S (.DIODE(_04248_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07659__A (.DIODE(_04248_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout286_A (.DIODE(_04249_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout284_A (.DIODE(_04249_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout283_A (.DIODE(_04249_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout282_A (.DIODE(_04249_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout267_A (.DIODE(_04251_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout265_A (.DIODE(_04251_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07781__S (.DIODE(_04251_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07771__S (.DIODE(_04251_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08932__A2 (.DIODE(_04254_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08927__A2 (.DIODE(_04254_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08926__A (.DIODE(_04254_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08908__A2_N (.DIODE(_04254_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07664__B (.DIODE(_04254_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09190__A2 (.DIODE(_04255_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09057__B (.DIODE(_04255_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08929__B (.DIODE(_04255_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08923__S (.DIODE(_04255_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08920__S (.DIODE(_04255_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08916__S (.DIODE(_04255_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08907__B (.DIODE(_04255_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08719__A2 (.DIODE(_04255_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07763__B (.DIODE(_04255_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07665__B (.DIODE(_04255_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout263_A (.DIODE(_04256_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout261_A (.DIODE(_04256_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout260_A (.DIODE(_04256_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout259_A (.DIODE(_04256_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09313__A (.DIODE(_04257_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09191__A2 (.DIODE(_04257_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09059__B (.DIODE(_04257_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09058__B (.DIODE(_04257_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07997__A2 (.DIODE(_04257_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07994__B1 (.DIODE(_04257_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07718__B1 (.DIODE(_04257_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07714__A1 (.DIODE(_04257_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07675__B1 (.DIODE(_04257_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07671__B1 (.DIODE(_04257_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout386_A (.DIODE(_04612_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout374_A (.DIODE(_04612_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout370_A (.DIODE(_04612_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout206_A (.DIODE(_04615_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout195_A (.DIODE(_04615_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout192_A (.DIODE(_04615_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout189_A (.DIODE(_04616_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout177_A (.DIODE(_04616_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout174_A (.DIODE(_04616_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08430__S (.DIODE(_04772_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08428__S (.DIODE(_04772_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08426__S (.DIODE(_04772_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08424__S (.DIODE(_04772_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08422__S (.DIODE(_04772_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08420__S (.DIODE(_04772_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08418__S (.DIODE(_04772_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08416__S (.DIODE(_04772_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08691__A2 (.DIODE(_04861_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08667__B2 (.DIODE(_04861_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08642__B (.DIODE(_04861_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08667__A2 (.DIODE(_04866_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08663__B (.DIODE(_04866_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08660__B1_N (.DIODE(_04866_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08658__A (.DIODE(_04866_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08655__B1 (.DIODE(_04866_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08653__A3 (.DIODE(_04866_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08650__B (.DIODE(_04866_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08649__B1 (.DIODE(_04866_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08666__B1 (.DIODE(_04868_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08665__A2 (.DIODE(_04868_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08662__B2 (.DIODE(_04868_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08657__B2 (.DIODE(_04868_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08651__B (.DIODE(_04868_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout325_A (.DIODE(_04917_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout324_A (.DIODE(_04917_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout323_A (.DIODE(_04917_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08776__B1 (.DIODE(_04917_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08934__B (.DIODE(_05059_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08933__A2 (.DIODE(_05059_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08932__B1 (.DIODE(_05059_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08931__S (.DIODE(_05059_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08928__S (.DIODE(_05059_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08924__S (.DIODE(_05059_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08921__S (.DIODE(_05059_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08917__S (.DIODE(_05059_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout322_A (.DIODE(_05075_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08936__A (.DIODE(_05075_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout227_A (.DIODE(_05253_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout223_A (.DIODE(_05253_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(en),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(gpio_in[10]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(gpio_in[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(gpio_in[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(gpio_in[4]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(gpio_in[5]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(gpio_in[6]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(gpio_in[7]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(gpio_in[8]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(gpio_in[9]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(nrst),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08031__A (.DIODE(\top.CB_read_complete ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08030__A (.DIODE(\top.CB_read_complete ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05964__A1 (.DIODE(\top.CB_read_complete ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05496__A (.DIODE(\top.CB_read_complete ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05495__A (.DIODE(\top.CB_read_complete ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09055__A1 (.DIODE(\top.CB_write_complete ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08036__B (.DIODE(\top.CB_write_complete ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08029__A (.DIODE(\top.CB_write_complete ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05965__B1 (.DIODE(\top.CB_write_complete ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05496__B (.DIODE(\top.CB_write_complete ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05495__B (.DIODE(\top.CB_write_complete ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09017__B2 (.DIODE(\top.TRN_char_index[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08837__C (.DIODE(\top.TRN_char_index[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06349__S (.DIODE(\top.TRN_char_index[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06325__B (.DIODE(\top.TRN_char_index[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06178__B (.DIODE(\top.TRN_char_index[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05738__A0 (.DIODE(\top.TRN_char_index[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09050__A0 (.DIODE(\top.WB.CPU_DAT_O[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08968__A0 (.DIODE(\top.WB.CPU_DAT_O[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08902__A1 (.DIODE(\top.WB.CPU_DAT_O[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06001__A0 (.DIODE(\top.WB.CPU_DAT_O[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05961__B2 (.DIODE(\top.WB.CPU_DAT_O[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05898__A1 (.DIODE(\top.WB.CPU_DAT_O[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05776__B2 (.DIODE(\top.WB.CPU_DAT_O[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05486__B2 (.DIODE(\top.WB.CPU_DAT_O[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09040__A0 (.DIODE(\top.WB.CPU_DAT_O[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08958__A0 (.DIODE(\top.WB.CPU_DAT_O[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08892__A1 (.DIODE(\top.WB.CPU_DAT_O[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05991__A0 (.DIODE(\top.WB.CPU_DAT_O[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05951__B2 (.DIODE(\top.WB.CPU_DAT_O[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05888__A1 (.DIODE(\top.WB.CPU_DAT_O[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05766__B2 (.DIODE(\top.WB.CPU_DAT_O[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05476__B2 (.DIODE(\top.WB.CPU_DAT_O[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09039__A0 (.DIODE(\top.WB.CPU_DAT_O[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08957__A0 (.DIODE(\top.WB.CPU_DAT_O[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08891__A1 (.DIODE(\top.WB.CPU_DAT_O[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05990__A0 (.DIODE(\top.WB.CPU_DAT_O[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05950__B2 (.DIODE(\top.WB.CPU_DAT_O[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05887__A1 (.DIODE(\top.WB.CPU_DAT_O[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05765__B2 (.DIODE(\top.WB.CPU_DAT_O[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05475__B2 (.DIODE(\top.WB.CPU_DAT_O[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09038__A0 (.DIODE(\top.WB.CPU_DAT_O[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08956__A0 (.DIODE(\top.WB.CPU_DAT_O[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08890__A1 (.DIODE(\top.WB.CPU_DAT_O[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05989__A0 (.DIODE(\top.WB.CPU_DAT_O[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05949__B2 (.DIODE(\top.WB.CPU_DAT_O[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05886__A1 (.DIODE(\top.WB.CPU_DAT_O[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05764__B2 (.DIODE(\top.WB.CPU_DAT_O[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05474__B2 (.DIODE(\top.WB.CPU_DAT_O[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09037__A0 (.DIODE(\top.WB.CPU_DAT_O[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08955__A0 (.DIODE(\top.WB.CPU_DAT_O[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08889__A1 (.DIODE(\top.WB.CPU_DAT_O[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05988__A0 (.DIODE(\top.WB.CPU_DAT_O[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05948__B2 (.DIODE(\top.WB.CPU_DAT_O[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05885__A1 (.DIODE(\top.WB.CPU_DAT_O[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05763__B2 (.DIODE(\top.WB.CPU_DAT_O[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05473__B2 (.DIODE(\top.WB.CPU_DAT_O[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09036__A0 (.DIODE(\top.WB.CPU_DAT_O[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09006__A0 (.DIODE(\top.WB.CPU_DAT_O[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08987__A0 (.DIODE(\top.WB.CPU_DAT_O[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08954__A0 (.DIODE(\top.WB.CPU_DAT_O[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08888__A1 (.DIODE(\top.WB.CPU_DAT_O[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05987__A0 (.DIODE(\top.WB.CPU_DAT_O[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05947__B2 (.DIODE(\top.WB.CPU_DAT_O[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05884__A1 (.DIODE(\top.WB.CPU_DAT_O[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05472__B2 (.DIODE(\top.WB.CPU_DAT_O[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09035__A0 (.DIODE(\top.WB.CPU_DAT_O[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09005__A0 (.DIODE(\top.WB.CPU_DAT_O[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08986__A0 (.DIODE(\top.WB.CPU_DAT_O[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08953__A0 (.DIODE(\top.WB.CPU_DAT_O[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08887__A1 (.DIODE(\top.WB.CPU_DAT_O[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05986__A0 (.DIODE(\top.WB.CPU_DAT_O[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05946__B2 (.DIODE(\top.WB.CPU_DAT_O[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05883__A1 (.DIODE(\top.WB.CPU_DAT_O[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05471__B2 (.DIODE(\top.WB.CPU_DAT_O[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09034__A0 (.DIODE(\top.WB.CPU_DAT_O[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09004__A0 (.DIODE(\top.WB.CPU_DAT_O[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08985__A0 (.DIODE(\top.WB.CPU_DAT_O[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08952__A0 (.DIODE(\top.WB.CPU_DAT_O[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08886__A1 (.DIODE(\top.WB.CPU_DAT_O[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05985__A0 (.DIODE(\top.WB.CPU_DAT_O[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05945__B2 (.DIODE(\top.WB.CPU_DAT_O[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05882__A1 (.DIODE(\top.WB.CPU_DAT_O[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05470__B2 (.DIODE(\top.WB.CPU_DAT_O[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09033__A0 (.DIODE(\top.WB.CPU_DAT_O[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09003__A0 (.DIODE(\top.WB.CPU_DAT_O[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08984__A0 (.DIODE(\top.WB.CPU_DAT_O[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08951__A0 (.DIODE(\top.WB.CPU_DAT_O[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08885__A1 (.DIODE(\top.WB.CPU_DAT_O[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05984__A0 (.DIODE(\top.WB.CPU_DAT_O[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05944__B2 (.DIODE(\top.WB.CPU_DAT_O[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05881__A1 (.DIODE(\top.WB.CPU_DAT_O[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05469__B2 (.DIODE(\top.WB.CPU_DAT_O[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09032__A0 (.DIODE(\top.WB.CPU_DAT_O[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09002__A0 (.DIODE(\top.WB.CPU_DAT_O[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08983__A0 (.DIODE(\top.WB.CPU_DAT_O[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08950__A0 (.DIODE(\top.WB.CPU_DAT_O[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08884__A1 (.DIODE(\top.WB.CPU_DAT_O[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05983__A0 (.DIODE(\top.WB.CPU_DAT_O[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05943__B2 (.DIODE(\top.WB.CPU_DAT_O[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05880__A1 (.DIODE(\top.WB.CPU_DAT_O[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05468__B2 (.DIODE(\top.WB.CPU_DAT_O[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09031__A0 (.DIODE(\top.WB.CPU_DAT_O[19] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09001__A0 (.DIODE(\top.WB.CPU_DAT_O[19] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08982__A0 (.DIODE(\top.WB.CPU_DAT_O[19] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08949__A0 (.DIODE(\top.WB.CPU_DAT_O[19] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08883__A1 (.DIODE(\top.WB.CPU_DAT_O[19] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05982__A0 (.DIODE(\top.WB.CPU_DAT_O[19] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05942__B2 (.DIODE(\top.WB.CPU_DAT_O[19] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05879__A1 (.DIODE(\top.WB.CPU_DAT_O[19] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05467__B2 (.DIODE(\top.WB.CPU_DAT_O[19] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09049__A0 (.DIODE(\top.WB.CPU_DAT_O[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08967__A0 (.DIODE(\top.WB.CPU_DAT_O[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08901__A1 (.DIODE(\top.WB.CPU_DAT_O[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06000__A0 (.DIODE(\top.WB.CPU_DAT_O[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05960__B2 (.DIODE(\top.WB.CPU_DAT_O[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05897__A1 (.DIODE(\top.WB.CPU_DAT_O[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05775__B2 (.DIODE(\top.WB.CPU_DAT_O[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05485__B2 (.DIODE(\top.WB.CPU_DAT_O[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09030__A0 (.DIODE(\top.WB.CPU_DAT_O[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09000__A0 (.DIODE(\top.WB.CPU_DAT_O[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08981__A0 (.DIODE(\top.WB.CPU_DAT_O[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08948__A0 (.DIODE(\top.WB.CPU_DAT_O[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08882__A1 (.DIODE(\top.WB.CPU_DAT_O[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05981__A0 (.DIODE(\top.WB.CPU_DAT_O[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05941__B2 (.DIODE(\top.WB.CPU_DAT_O[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05878__A1 (.DIODE(\top.WB.CPU_DAT_O[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05466__B2 (.DIODE(\top.WB.CPU_DAT_O[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09029__A0 (.DIODE(\top.WB.CPU_DAT_O[21] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08999__A0 (.DIODE(\top.WB.CPU_DAT_O[21] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08980__A0 (.DIODE(\top.WB.CPU_DAT_O[21] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08947__A0 (.DIODE(\top.WB.CPU_DAT_O[21] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08881__A1 (.DIODE(\top.WB.CPU_DAT_O[21] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05980__A0 (.DIODE(\top.WB.CPU_DAT_O[21] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05940__B2 (.DIODE(\top.WB.CPU_DAT_O[21] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05877__A1 (.DIODE(\top.WB.CPU_DAT_O[21] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05465__B2 (.DIODE(\top.WB.CPU_DAT_O[21] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09028__A0 (.DIODE(\top.WB.CPU_DAT_O[22] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08998__A0 (.DIODE(\top.WB.CPU_DAT_O[22] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08979__A0 (.DIODE(\top.WB.CPU_DAT_O[22] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08946__A0 (.DIODE(\top.WB.CPU_DAT_O[22] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08880__A1 (.DIODE(\top.WB.CPU_DAT_O[22] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05979__A0 (.DIODE(\top.WB.CPU_DAT_O[22] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05939__B2 (.DIODE(\top.WB.CPU_DAT_O[22] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05876__A1 (.DIODE(\top.WB.CPU_DAT_O[22] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05464__B2 (.DIODE(\top.WB.CPU_DAT_O[22] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09027__A0 (.DIODE(\top.WB.CPU_DAT_O[23] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08997__A0 (.DIODE(\top.WB.CPU_DAT_O[23] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08978__A0 (.DIODE(\top.WB.CPU_DAT_O[23] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08945__A0 (.DIODE(\top.WB.CPU_DAT_O[23] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08879__A1 (.DIODE(\top.WB.CPU_DAT_O[23] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05978__A0 (.DIODE(\top.WB.CPU_DAT_O[23] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05938__B2 (.DIODE(\top.WB.CPU_DAT_O[23] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05875__A1 (.DIODE(\top.WB.CPU_DAT_O[23] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05463__B2 (.DIODE(\top.WB.CPU_DAT_O[23] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09026__A0 (.DIODE(\top.WB.CPU_DAT_O[24] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08996__A0 (.DIODE(\top.WB.CPU_DAT_O[24] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08977__A0 (.DIODE(\top.WB.CPU_DAT_O[24] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08944__A0 (.DIODE(\top.WB.CPU_DAT_O[24] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08878__A1 (.DIODE(\top.WB.CPU_DAT_O[24] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05977__A0 (.DIODE(\top.WB.CPU_DAT_O[24] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05937__B2 (.DIODE(\top.WB.CPU_DAT_O[24] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05874__A1 (.DIODE(\top.WB.CPU_DAT_O[24] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05462__B2 (.DIODE(\top.WB.CPU_DAT_O[24] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09025__A0 (.DIODE(\top.WB.CPU_DAT_O[25] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08995__A0 (.DIODE(\top.WB.CPU_DAT_O[25] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08976__A0 (.DIODE(\top.WB.CPU_DAT_O[25] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08943__A0 (.DIODE(\top.WB.CPU_DAT_O[25] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08877__A1 (.DIODE(\top.WB.CPU_DAT_O[25] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05976__A0 (.DIODE(\top.WB.CPU_DAT_O[25] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05936__B2 (.DIODE(\top.WB.CPU_DAT_O[25] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05873__A1 (.DIODE(\top.WB.CPU_DAT_O[25] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05461__B2 (.DIODE(\top.WB.CPU_DAT_O[25] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09024__A0 (.DIODE(\top.WB.CPU_DAT_O[26] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08994__A0 (.DIODE(\top.WB.CPU_DAT_O[26] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08975__A0 (.DIODE(\top.WB.CPU_DAT_O[26] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08942__A0 (.DIODE(\top.WB.CPU_DAT_O[26] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08876__A1 (.DIODE(\top.WB.CPU_DAT_O[26] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05975__A0 (.DIODE(\top.WB.CPU_DAT_O[26] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05935__B2 (.DIODE(\top.WB.CPU_DAT_O[26] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05872__A1 (.DIODE(\top.WB.CPU_DAT_O[26] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05460__B2 (.DIODE(\top.WB.CPU_DAT_O[26] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09023__A0 (.DIODE(\top.WB.CPU_DAT_O[27] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08993__A0 (.DIODE(\top.WB.CPU_DAT_O[27] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08974__A0 (.DIODE(\top.WB.CPU_DAT_O[27] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08941__A0 (.DIODE(\top.WB.CPU_DAT_O[27] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08875__A1 (.DIODE(\top.WB.CPU_DAT_O[27] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05974__A0 (.DIODE(\top.WB.CPU_DAT_O[27] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05934__B2 (.DIODE(\top.WB.CPU_DAT_O[27] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05871__A1 (.DIODE(\top.WB.CPU_DAT_O[27] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05459__B2 (.DIODE(\top.WB.CPU_DAT_O[27] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09022__A0 (.DIODE(\top.WB.CPU_DAT_O[28] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08992__A0 (.DIODE(\top.WB.CPU_DAT_O[28] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08973__A0 (.DIODE(\top.WB.CPU_DAT_O[28] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08940__A0 (.DIODE(\top.WB.CPU_DAT_O[28] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08874__A1 (.DIODE(\top.WB.CPU_DAT_O[28] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05973__A0 (.DIODE(\top.WB.CPU_DAT_O[28] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05933__B2 (.DIODE(\top.WB.CPU_DAT_O[28] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05870__A1 (.DIODE(\top.WB.CPU_DAT_O[28] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05458__B2 (.DIODE(\top.WB.CPU_DAT_O[28] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09021__A0 (.DIODE(\top.WB.CPU_DAT_O[29] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08991__A0 (.DIODE(\top.WB.CPU_DAT_O[29] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08972__A0 (.DIODE(\top.WB.CPU_DAT_O[29] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08939__A0 (.DIODE(\top.WB.CPU_DAT_O[29] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08873__A1 (.DIODE(\top.WB.CPU_DAT_O[29] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05972__A0 (.DIODE(\top.WB.CPU_DAT_O[29] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05932__B2 (.DIODE(\top.WB.CPU_DAT_O[29] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05869__A1 (.DIODE(\top.WB.CPU_DAT_O[29] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05457__B2 (.DIODE(\top.WB.CPU_DAT_O[29] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09048__A0 (.DIODE(\top.WB.CPU_DAT_O[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08966__A0 (.DIODE(\top.WB.CPU_DAT_O[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08900__A1 (.DIODE(\top.WB.CPU_DAT_O[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05999__A0 (.DIODE(\top.WB.CPU_DAT_O[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05959__B2 (.DIODE(\top.WB.CPU_DAT_O[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05896__A1 (.DIODE(\top.WB.CPU_DAT_O[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05774__B2 (.DIODE(\top.WB.CPU_DAT_O[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05484__B2 (.DIODE(\top.WB.CPU_DAT_O[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09020__A0 (.DIODE(\top.WB.CPU_DAT_O[30] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08990__A0 (.DIODE(\top.WB.CPU_DAT_O[30] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08971__A0 (.DIODE(\top.WB.CPU_DAT_O[30] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08938__A0 (.DIODE(\top.WB.CPU_DAT_O[30] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08872__A1 (.DIODE(\top.WB.CPU_DAT_O[30] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05971__A0 (.DIODE(\top.WB.CPU_DAT_O[30] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05931__B2 (.DIODE(\top.WB.CPU_DAT_O[30] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05868__A1 (.DIODE(\top.WB.CPU_DAT_O[30] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05456__B2 (.DIODE(\top.WB.CPU_DAT_O[30] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09019__A0 (.DIODE(\top.WB.CPU_DAT_O[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08989__A0 (.DIODE(\top.WB.CPU_DAT_O[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08970__A0 (.DIODE(\top.WB.CPU_DAT_O[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08937__A0 (.DIODE(\top.WB.CPU_DAT_O[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08871__A1 (.DIODE(\top.WB.CPU_DAT_O[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05970__A0 (.DIODE(\top.WB.CPU_DAT_O[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05930__B2 (.DIODE(\top.WB.CPU_DAT_O[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05867__A1 (.DIODE(\top.WB.CPU_DAT_O[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05455__B2 (.DIODE(\top.WB.CPU_DAT_O[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09047__A0 (.DIODE(\top.WB.CPU_DAT_O[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08965__A0 (.DIODE(\top.WB.CPU_DAT_O[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08899__A1 (.DIODE(\top.WB.CPU_DAT_O[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05998__A0 (.DIODE(\top.WB.CPU_DAT_O[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05958__B2 (.DIODE(\top.WB.CPU_DAT_O[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05895__A1 (.DIODE(\top.WB.CPU_DAT_O[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05773__B2 (.DIODE(\top.WB.CPU_DAT_O[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05483__B2 (.DIODE(\top.WB.CPU_DAT_O[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09046__A0 (.DIODE(\top.WB.CPU_DAT_O[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08964__A0 (.DIODE(\top.WB.CPU_DAT_O[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08898__A1 (.DIODE(\top.WB.CPU_DAT_O[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05997__A0 (.DIODE(\top.WB.CPU_DAT_O[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05957__B2 (.DIODE(\top.WB.CPU_DAT_O[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05894__A1 (.DIODE(\top.WB.CPU_DAT_O[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05772__B2 (.DIODE(\top.WB.CPU_DAT_O[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05482__B2 (.DIODE(\top.WB.CPU_DAT_O[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09045__A0 (.DIODE(\top.WB.CPU_DAT_O[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08963__A0 (.DIODE(\top.WB.CPU_DAT_O[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08897__A1 (.DIODE(\top.WB.CPU_DAT_O[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05996__A0 (.DIODE(\top.WB.CPU_DAT_O[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05956__B2 (.DIODE(\top.WB.CPU_DAT_O[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05893__A1 (.DIODE(\top.WB.CPU_DAT_O[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05771__B2 (.DIODE(\top.WB.CPU_DAT_O[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05481__B2 (.DIODE(\top.WB.CPU_DAT_O[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09044__A0 (.DIODE(\top.WB.CPU_DAT_O[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08962__A0 (.DIODE(\top.WB.CPU_DAT_O[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08896__A1 (.DIODE(\top.WB.CPU_DAT_O[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05995__A0 (.DIODE(\top.WB.CPU_DAT_O[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05955__B2 (.DIODE(\top.WB.CPU_DAT_O[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05892__A1 (.DIODE(\top.WB.CPU_DAT_O[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05770__B2 (.DIODE(\top.WB.CPU_DAT_O[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05480__B2 (.DIODE(\top.WB.CPU_DAT_O[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09043__A0 (.DIODE(\top.WB.CPU_DAT_O[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08961__A0 (.DIODE(\top.WB.CPU_DAT_O[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08895__A1 (.DIODE(\top.WB.CPU_DAT_O[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05994__A0 (.DIODE(\top.WB.CPU_DAT_O[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05954__B2 (.DIODE(\top.WB.CPU_DAT_O[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05891__A1 (.DIODE(\top.WB.CPU_DAT_O[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05769__B2 (.DIODE(\top.WB.CPU_DAT_O[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05479__B2 (.DIODE(\top.WB.CPU_DAT_O[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09042__A0 (.DIODE(\top.WB.CPU_DAT_O[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08960__A0 (.DIODE(\top.WB.CPU_DAT_O[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08894__A1 (.DIODE(\top.WB.CPU_DAT_O[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05993__A0 (.DIODE(\top.WB.CPU_DAT_O[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05953__B2 (.DIODE(\top.WB.CPU_DAT_O[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05890__A1 (.DIODE(\top.WB.CPU_DAT_O[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05768__B2 (.DIODE(\top.WB.CPU_DAT_O[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05478__B2 (.DIODE(\top.WB.CPU_DAT_O[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09041__A0 (.DIODE(\top.WB.CPU_DAT_O[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08959__A0 (.DIODE(\top.WB.CPU_DAT_O[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08893__A1 (.DIODE(\top.WB.CPU_DAT_O[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05992__A0 (.DIODE(\top.WB.CPU_DAT_O[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05952__B2 (.DIODE(\top.WB.CPU_DAT_O[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05889__A1 (.DIODE(\top.WB.CPU_DAT_O[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05767__B2 (.DIODE(\top.WB.CPU_DAT_O[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05477__B2 (.DIODE(\top.WB.CPU_DAT_O[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09175__A1 (.DIODE(\top.WB.curr_state[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05487__B (.DIODE(\top.WB.curr_state[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05452__A (.DIODE(\top.WB.curr_state[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05451__A (.DIODE(\top.WB.curr_state[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06041__C_N (.DIODE(\top.WB.prev_BUSY_O ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05860__B (.DIODE(\top.WB.prev_BUSY_O ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05454__C_N (.DIODE(\top.WB.prev_BUSY_O ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05453__B (.DIODE(\top.WB.prev_BUSY_O ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09233__A1 (.DIODE(\top.cb_syn.char_index[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08420__A0 (.DIODE(\top.cb_syn.char_index[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06239__A (.DIODE(\top.cb_syn.char_index[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06238__A1 (.DIODE(\top.cb_syn.char_index[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06172__A (.DIODE(\top.cb_syn.char_index[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06166__A2 (.DIODE(\top.cb_syn.char_index[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06161__A (.DIODE(\top.cb_syn.char_index[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout520_A (.DIODE(\top.cb_syn.char_path_n[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08660__A1 (.DIODE(\top.cb_syn.char_path_n[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05421__A (.DIODE(\top.cb_syn.char_path_n[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08559__A1 (.DIODE(\top.cb_syn.char_path_n[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09194__A1 (.DIODE(\top.cb_syn.char_path_n[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09166__A_N (.DIODE(\top.cb_syn.char_path_n[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09054__A1 (.DIODE(\top.cb_syn.char_path_n[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08619__A0 (.DIODE(\top.cb_syn.char_path_n[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08558__A1 (.DIODE(\top.cb_syn.char_path_n[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08406__A1 (.DIODE(\top.cb_syn.char_path_n[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08403__B2 (.DIODE(\top.cb_syn.char_path_n[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08051__A (.DIODE(\top.cb_syn.char_path_n[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07548__A1 (.DIODE(\top.cb_syn.char_path_n[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09158__A_N (.DIODE(\top.cb_syn.char_path_n[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08619__A1 (.DIODE(\top.cb_syn.char_path_n[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08557__A1 (.DIODE(\top.cb_syn.char_path_n[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08405__A1 (.DIODE(\top.cb_syn.char_path_n[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08404__A1 (.DIODE(\top.cb_syn.char_path_n[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08401__B2 (.DIODE(\top.cb_syn.char_path_n[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08052__A (.DIODE(\top.cb_syn.char_path_n[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07548__A0 (.DIODE(\top.cb_syn.char_path_n[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08608__A3 (.DIODE(\top.cb_syn.char_path_n[32] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08527__A1 (.DIODE(\top.cb_syn.char_path_n[32] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08345__A1 (.DIODE(\top.cb_syn.char_path_n[32] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08344__A1 (.DIODE(\top.cb_syn.char_path_n[32] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08341__B2 (.DIODE(\top.cb_syn.char_path_n[32] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07551__A2 (.DIODE(\top.cb_syn.char_path_n[32] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08635__A0 (.DIODE(\top.cb_syn.char_path_n[33] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08526__A1 (.DIODE(\top.cb_syn.char_path_n[33] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08343__A1 (.DIODE(\top.cb_syn.char_path_n[33] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08342__A1 (.DIODE(\top.cb_syn.char_path_n[33] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08339__B2 (.DIODE(\top.cb_syn.char_path_n[33] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07563__A1 (.DIODE(\top.cb_syn.char_path_n[33] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08585__A0 (.DIODE(\top.cb_syn.char_path_n[65] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08494__A1 (.DIODE(\top.cb_syn.char_path_n[65] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08279__A1 (.DIODE(\top.cb_syn.char_path_n[65] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08278__A1 (.DIODE(\top.cb_syn.char_path_n[65] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08275__B2 (.DIODE(\top.cb_syn.char_path_n[65] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07532__A1 (.DIODE(\top.cb_syn.char_path_n[65] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08620__A2 (.DIODE(\top.cb_syn.char_path_n[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08552__A1 (.DIODE(\top.cb_syn.char_path_n[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08395__A1 (.DIODE(\top.cb_syn.char_path_n[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08394__A1 (.DIODE(\top.cb_syn.char_path_n[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08391__B2 (.DIODE(\top.cb_syn.char_path_n[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07547__A3 (.DIODE(\top.cb_syn.char_path_n[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08574__A3 (.DIODE(\top.cb_syn.char_path_n[88] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08471__A1 (.DIODE(\top.cb_syn.char_path_n[88] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08233__A1 (.DIODE(\top.cb_syn.char_path_n[88] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08232__A1 (.DIODE(\top.cb_syn.char_path_n[88] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08229__B2 (.DIODE(\top.cb_syn.char_path_n[88] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07538__A2 (.DIODE(\top.cb_syn.char_path_n[88] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08620__A3 (.DIODE(\top.cb_syn.char_path_n[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08551__A1 (.DIODE(\top.cb_syn.char_path_n[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08393__A1 (.DIODE(\top.cb_syn.char_path_n[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08392__A1 (.DIODE(\top.cb_syn.char_path_n[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08389__B2 (.DIODE(\top.cb_syn.char_path_n[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07547__A2 (.DIODE(\top.cb_syn.char_path_n[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08578__A3 (.DIODE(\top.cb_syn.char_path_n[96] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08463__A1 (.DIODE(\top.cb_syn.char_path_n[96] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08217__A1 (.DIODE(\top.cb_syn.char_path_n[96] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08216__A1 (.DIODE(\top.cb_syn.char_path_n[96] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08213__B2 (.DIODE(\top.cb_syn.char_path_n[96] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07535__A2 (.DIODE(\top.cb_syn.char_path_n[96] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08594__A0 (.DIODE(\top.cb_syn.char_path_n[97] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08462__A1 (.DIODE(\top.cb_syn.char_path_n[97] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08215__A1 (.DIODE(\top.cb_syn.char_path_n[97] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08214__A1 (.DIODE(\top.cb_syn.char_path_n[97] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08211__B2 (.DIODE(\top.cb_syn.char_path_n[97] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07517__A1 (.DIODE(\top.cb_syn.char_path_n[97] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08594__A1 (.DIODE(\top.cb_syn.char_path_n[98] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08461__A1 (.DIODE(\top.cb_syn.char_path_n[98] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08213__A1 (.DIODE(\top.cb_syn.char_path_n[98] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08212__A1 (.DIODE(\top.cb_syn.char_path_n[98] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08209__B2 (.DIODE(\top.cb_syn.char_path_n[98] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07517__A0 (.DIODE(\top.cb_syn.char_path_n[98] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08659__A1 (.DIODE(\top.cb_syn.end_cnt[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08638__A1 (.DIODE(\top.cb_syn.end_cnt[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08622__A (.DIODE(\top.cb_syn.end_cnt[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08614__A1 (.DIODE(\top.cb_syn.end_cnt[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08604__B1 (.DIODE(\top.cb_syn.end_cnt[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08597__B2 (.DIODE(\top.cb_syn.end_cnt[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08588__B2 (.DIODE(\top.cb_syn.end_cnt[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08580__A1 (.DIODE(\top.cb_syn.end_cnt[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08570__A (.DIODE(\top.cb_syn.end_cnt[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05424__A (.DIODE(\top.cb_syn.end_cnt[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08652__S (.DIODE(\top.cb_syn.end_cnt[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08641__A1 (.DIODE(\top.cb_syn.end_cnt[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08640__B1 (.DIODE(\top.cb_syn.end_cnt[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08572__B2 (.DIODE(\top.cb_syn.end_cnt[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06947__B2 (.DIODE(\top.compVal[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06887__A0 (.DIODE(\top.compVal[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06731__B2 (.DIODE(\top.compVal[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06598__B (.DIODE(\top.compVal[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05951__A1 (.DIODE(\top.compVal[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05319__A (.DIODE(\top.compVal[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09201__B (.DIODE(\top.controller.fin_reg[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09199__B (.DIODE(\top.controller.fin_reg[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09196__D_N (.DIODE(\top.controller.fin_reg[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09178__B (.DIODE(\top.controller.fin_reg[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout469_A (.DIODE(\top.controller.state_reg[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout466_A (.DIODE(\top.controller.state_reg[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout454_A (.DIODE(\top.controller.state_reg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06365__C1 (.DIODE(\top.controller.state_reg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06011__B (.DIODE(\top.controller.state_reg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout452_A (.DIODE(\top.controller.state_reg[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06309__C1 (.DIODE(\top.controller.state_reg[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06350__B2 (.DIODE(\top.controller.state_reg[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06125__B (.DIODE(\top.controller.state_reg[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07426__B2 (.DIODE(\top.findLeastValue.histo_index[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07413__A0 (.DIODE(\top.findLeastValue.histo_index[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07008__B2 (.DIODE(\top.findLeastValue.histo_index[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06996__B2 (.DIODE(\top.findLeastValue.histo_index[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06984__A1 (.DIODE(\top.findLeastValue.histo_index[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06336__B1 (.DIODE(\top.findLeastValue.histo_index[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06320__A1 (.DIODE(\top.findLeastValue.histo_index[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06318__A1 (.DIODE(\top.findLeastValue.histo_index[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06215__A (.DIODE(\top.findLeastValue.histo_index[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05488__D (.DIODE(\top.findLeastValue.histo_index[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07402__A0 (.DIODE(\top.findLeastValue.histo_index[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06976__A1 (.DIODE(\top.findLeastValue.histo_index[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06973__A1 (.DIODE(\top.findLeastValue.histo_index[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06162__B (.DIODE(\top.findLeastValue.histo_index[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05748__A1 (.DIODE(\top.findLeastValue.histo_index[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05743__B (.DIODE(\top.findLeastValue.histo_index[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05742__B (.DIODE(\top.findLeastValue.histo_index[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05490__A (.DIODE(\top.findLeastValue.histo_index[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05384__A (.DIODE(\top.findLeastValue.histo_index[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08011__A1 (.DIODE(\top.findLeastValue.least1[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07708__A1 (.DIODE(\top.findLeastValue.least1[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07707__A1 (.DIODE(\top.findLeastValue.least1[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07428__A1 (.DIODE(\top.findLeastValue.least1[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07417__A1 (.DIODE(\top.findLeastValue.least1[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05807__D (.DIODE(\top.findLeastValue.least1[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08011__A0 (.DIODE(\top.findLeastValue.least2[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07756__A1 (.DIODE(\top.findLeastValue.least2[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07755__A1 (.DIODE(\top.findLeastValue.least2[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05811__D (.DIODE(\top.findLeastValue.least2[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05404__A (.DIODE(\top.findLeastValue.least2[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold773_A (.DIODE(\top.findLeastValue.sum[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07989__B2 (.DIODE(\top.findLeastValue.sum[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07986__A0 (.DIODE(\top.findLeastValue.sum[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07985__A1 (.DIODE(\top.findLeastValue.sum[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07934__B2 (.DIODE(\top.findLeastValue.sum[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07931__A1 (.DIODE(\top.findLeastValue.sum[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07930__A1 (.DIODE(\top.findLeastValue.sum[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07370__B2 (.DIODE(\top.findLeastValue.sum[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold608_A (.DIODE(\top.findLeastValue.sum[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07921__A1 (.DIODE(\top.findLeastValue.sum[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07920__A1 (.DIODE(\top.findLeastValue.sum[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07914__B2 (.DIODE(\top.findLeastValue.sum[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07911__A0 (.DIODE(\top.findLeastValue.sum[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07910__A1 (.DIODE(\top.findLeastValue.sum[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07358__B2 (.DIODE(\top.findLeastValue.sum[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold798_A (.DIODE(\top.findLeastValue.sum[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07984__B2 (.DIODE(\top.findLeastValue.sum[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07981__A1 (.DIODE(\top.findLeastValue.sum[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07980__A1 (.DIODE(\top.findLeastValue.sum[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07979__B2 (.DIODE(\top.findLeastValue.sum[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07976__A0 (.DIODE(\top.findLeastValue.sum[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07975__A1 (.DIODE(\top.findLeastValue.sum[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07395__B2 (.DIODE(\top.findLeastValue.sum[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold764_A (.DIODE(\top.findLeastValue.sum[33] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07824__B2 (.DIODE(\top.findLeastValue.sum[33] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07821__A1 (.DIODE(\top.findLeastValue.sum[33] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07820__A1 (.DIODE(\top.findLeastValue.sum[33] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07819__B2 (.DIODE(\top.findLeastValue.sum[34] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07816__A0 (.DIODE(\top.findLeastValue.sum[34] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07815__A1 (.DIODE(\top.findLeastValue.sum[34] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07286__B2 (.DIODE(\top.findLeastValue.sum[34] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07814__B2 (.DIODE(\top.findLeastValue.sum[35] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07811__A0 (.DIODE(\top.findLeastValue.sum[35] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07810__A1 (.DIODE(\top.findLeastValue.sum[35] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07284__B2 (.DIODE(\top.findLeastValue.sum[35] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold745_A (.DIODE(\top.findLeastValue.sum[37] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07804__B2 (.DIODE(\top.findLeastValue.sum[37] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07801__A1 (.DIODE(\top.findLeastValue.sum[37] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07800__A1 (.DIODE(\top.findLeastValue.sum[37] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07799__B2 (.DIODE(\top.findLeastValue.sum[38] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07796__A1 (.DIODE(\top.findLeastValue.sum[38] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07795__A1 (.DIODE(\top.findLeastValue.sum[38] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07271__A1 (.DIODE(\top.findLeastValue.sum[38] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold732_A (.DIODE(\top.findLeastValue.sum[39] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07794__B2 (.DIODE(\top.findLeastValue.sum[39] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07791__A1 (.DIODE(\top.findLeastValue.sum[39] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07790__A1 (.DIODE(\top.findLeastValue.sum[39] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold840_A (.DIODE(\top.findLeastValue.sum[41] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07784__B2 (.DIODE(\top.findLeastValue.sum[41] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07781__A1 (.DIODE(\top.findLeastValue.sum[41] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07780__A1 (.DIODE(\top.findLeastValue.sum[41] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold776_A (.DIODE(\top.findLeastValue.sum[43] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07774__B2 (.DIODE(\top.findLeastValue.sum[43] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07771__A1 (.DIODE(\top.findLeastValue.sum[43] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07770__A1 (.DIODE(\top.findLeastValue.sum[43] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07769__B2 (.DIODE(\top.findLeastValue.sum[44] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07766__A0 (.DIODE(\top.findLeastValue.sum[44] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07765__A1 (.DIODE(\top.findLeastValue.sum[44] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07249__B1 (.DIODE(\top.findLeastValue.sum[44] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold781_A (.DIODE(\top.findLeastValue.sum[45] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07764__B2 (.DIODE(\top.findLeastValue.sum[45] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07760__A1 (.DIODE(\top.findLeastValue.sum[45] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07759__A1 (.DIODE(\top.findLeastValue.sum[45] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07969__B2 (.DIODE(\top.findLeastValue.sum[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07966__A0 (.DIODE(\top.findLeastValue.sum[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07965__A1 (.DIODE(\top.findLeastValue.sum[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07391__B2 (.DIODE(\top.findLeastValue.sum[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07964__B2 (.DIODE(\top.findLeastValue.sum[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07961__A1 (.DIODE(\top.findLeastValue.sum[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07960__A1 (.DIODE(\top.findLeastValue.sum[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07389__B2 (.DIODE(\top.findLeastValue.sum[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07944__B2 (.DIODE(\top.findLeastValue.sum[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07941__A1 (.DIODE(\top.findLeastValue.sum[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07940__A1 (.DIODE(\top.findLeastValue.sum[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07376__B2 (.DIODE(\top.findLeastValue.sum[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07033__A (.DIODE(\top.findLeastValue.val1[46] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06911__A1 (.DIODE(\top.findLeastValue.val1[46] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06816__B2 (.DIODE(\top.findLeastValue.val1[46] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06686__B1 (.DIODE(\top.findLeastValue.val1[46] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold678_A (.DIODE(\top.hTree.node_reg[28] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05560__B2 (.DIODE(\top.hTree.node_reg[28] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold844_A (.DIODE(\top.hTree.node_reg[29] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05554__B2 (.DIODE(\top.hTree.node_reg[29] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09345__A1 (.DIODE(\top.hTree.node_reg[30] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05548__B2 (.DIODE(\top.hTree.node_reg[30] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09346__A1 (.DIODE(\top.hTree.node_reg[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05542__B2 (.DIODE(\top.hTree.node_reg[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold714_A (.DIODE(\top.hTree.node_reg[47] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05639__A1 (.DIODE(\top.hTree.node_reg[47] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold629_A (.DIODE(\top.hTree.node_reg[63] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05543__A1 (.DIODE(\top.hTree.node_reg[63] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09181__B1 (.DIODE(\top.hTree.write_HT_fin ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09084__B2 (.DIODE(\top.hTree.write_HT_fin ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08910__A (.DIODE(\top.hTree.write_HT_fin ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07663__A (.DIODE(\top.hTree.write_HT_fin ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07662__A (.DIODE(\top.hTree.write_HT_fin ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07658__A (.DIODE(\top.hTree.write_HT_fin ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06230__A1 (.DIODE(\top.hTree.write_HT_fin ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05865__B2 (.DIODE(\top.hTree.write_HT_fin ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05816__A (.DIODE(\top.hTree.write_HT_fin ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05301__A (.DIODE(\top.hTree.write_HT_fin ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09307__A1 (.DIODE(\top.header_synthesis.bit1 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06590__A1 (.DIODE(\top.header_synthesis.bit1 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09307__A3 (.DIODE(\top.header_synthesis.enable ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08842__A2 (.DIODE(\top.header_synthesis.enable ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08709__A1 (.DIODE(\top.header_synthesis.enable ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06572__A (.DIODE(\top.header_synthesis.enable ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05448__A (.DIODE(\top.header_synthesis.enable ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout549_A (.DIODE(\top.sram_interface.word_cnt[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout546_A (.DIODE(\top.sram_interface.word_cnt[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05581__A2 (.DIODE(\top.sram_interface.word_cnt[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05564__A2 (.DIODE(\top.sram_interface.word_cnt[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09144__B1 (.DIODE(\top.sram_interface.word_cnt[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09094__A2 (.DIODE(\top.sram_interface.word_cnt[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09084__A2 (.DIODE(\top.sram_interface.word_cnt[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09077__B1 (.DIODE(\top.sram_interface.word_cnt[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08969__B (.DIODE(\top.sram_interface.word_cnt[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05447__A (.DIODE(\top.sram_interface.word_cnt[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout541_A (.DIODE(\top.sram_interface.word_cnt[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout538_A (.DIODE(\top.sram_interface.word_cnt[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout537_A (.DIODE(\top.sram_interface.word_cnt[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout505_A (.DIODE(\top.translation.index[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08804__C1 (.DIODE(\top.translation.index[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08792__A1 (.DIODE(\top.translation.index[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08783__C1 (.DIODE(\top.translation.index[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09304__S (.DIODE(\top.translation.index[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08857__A1 (.DIODE(\top.translation.index[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08834__A1 (.DIODE(\top.translation.index[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08832__B1 (.DIODE(\top.translation.index[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05782__A (.DIODE(\top.translation.index[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08854__A (.DIODE(\top.translation.index[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08850__A1 (.DIODE(\top.translation.index[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08829__B1 (.DIODE(\top.translation.index[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08827__B1 (.DIODE(\top.translation.index[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08779__C1 (.DIODE(\top.translation.index[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08773__A1 (.DIODE(\top.translation.index[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05784__B (.DIODE(\top.translation.index[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05429__A (.DIODE(\top.translation.index[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08852__B2 (.DIODE(\top.translation.index[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08850__B1 (.DIODE(\top.translation.index[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08832__A1 (.DIODE(\top.translation.index[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08828__C1 (.DIODE(\top.translation.index[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08780__C1 (.DIODE(\top.translation.index[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05784__A (.DIODE(\top.translation.index[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05428__A (.DIODE(\top.translation.index[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05476__A1 (.DIODE(net3),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout877_A (.DIODE(net34),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout796_A (.DIODE(net34),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09307__A2 (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08842__B1 (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05778__C (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05777__B (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07492__A1 (.DIODE(net39),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05737__A1 (.DIODE(net39),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07487__A1 (.DIODE(net40),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05736__A1 (.DIODE(net40),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07482__A1 (.DIODE(net41),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05735__A1 (.DIODE(net41),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07476__A1 (.DIODE(net42),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05734__A1 (.DIODE(net42),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout712_A (.DIODE(net44),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout631_A (.DIODE(net44),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_output68_A (.DIODE(net68),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06313__A1 (.DIODE(net68),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout444_A (.DIODE(net72),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout441_A (.DIODE(net72),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05454__A (.DIODE(net72),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_output89_A (.DIODE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05586__A1 (.DIODE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_output93_A (.DIODE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05562__A1 (.DIODE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold826_A (.DIODE(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_output94_A (.DIODE(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold845_A (.DIODE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_output96_A (.DIODE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_output97_A (.DIODE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05544__A1 (.DIODE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06947__B1 (.DIODE(net113),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06948__B1 (.DIODE(net113),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06949__B1 (.DIODE(net113),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06913__B1 (.DIODE(net113),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06912__B1 (.DIODE(net113),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06946__B1 (.DIODE(net113),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06950__B1 (.DIODE(net113),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06951__B1 (.DIODE(net113),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06914__B1 (.DIODE(net113),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout112_A (.DIODE(net113),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout113_A (.DIODE(net114),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06922__B1 (.DIODE(net114),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06921__B1 (.DIODE(net114),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06920__B1 (.DIODE(net114),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06919__B1 (.DIODE(net114),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06924__B1 (.DIODE(net114),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06925__B1 (.DIODE(net114),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06923__B1 (.DIODE(net114),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06926__B1 (.DIODE(net114),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06929__B1 (.DIODE(net114),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06934__B1 (.DIODE(net115),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06933__B1 (.DIODE(net115),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06932__B1 (.DIODE(net115),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06931__B1 (.DIODE(net115),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06930__B1 (.DIODE(net115),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06928__B1 (.DIODE(net115),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06927__B1 (.DIODE(net115),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06938__B1 (.DIODE(net115),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06941__B1 (.DIODE(net115),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06940__B1 (.DIODE(net115),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06939__B1 (.DIODE(net116),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06944__B1 (.DIODE(net116),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06943__B1 (.DIODE(net116),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06942__B1 (.DIODE(net116),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06945__B1 (.DIODE(net116),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06936__B1 (.DIODE(net116),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06935__B1 (.DIODE(net116),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06937__B1 (.DIODE(net116),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout115_A (.DIODE(net116),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06858__B1 (.DIODE(net117),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06864__B1 (.DIODE(net117),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06862__B1 (.DIODE(net117),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06866__B1 (.DIODE(net117),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06868__B1 (.DIODE(net117),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06870__B1 (.DIODE(net117),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06856__B1 (.DIODE(net117),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06854__B1 (.DIODE(net117),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07404__B1 (.DIODE(net117),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07401__B1 (.DIODE(net117),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06848__B1 (.DIODE(net118),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06850__B1 (.DIODE(net118),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06842__B1 (.DIODE(net118),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06846__B1 (.DIODE(net118),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06852__B1 (.DIODE(net118),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06844__B1 (.DIODE(net118),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06840__B1 (.DIODE(net118),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06838__B1 (.DIODE(net118),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06836__B1 (.DIODE(net118),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06834__B1 (.DIODE(net118),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06820__B1 (.DIODE(net119),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06818__B1 (.DIODE(net119),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06816__B1 (.DIODE(net119),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06884__B1 (.DIODE(net119),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06822__B1 (.DIODE(net119),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06828__B1 (.DIODE(net119),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06826__B1 (.DIODE(net119),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06824__B1 (.DIODE(net119),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06830__B1 (.DIODE(net119),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06832__B1 (.DIODE(net119),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06894__B1 (.DIODE(net120),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06886__B1 (.DIODE(net120),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06882__B1 (.DIODE(net120),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06890__B1 (.DIODE(net120),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06904__B1 (.DIODE(net120),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06908__B1 (.DIODE(net120),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06906__B1 (.DIODE(net120),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06902__B1 (.DIODE(net120),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06898__B1 (.DIODE(net120),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06900__B1 (.DIODE(net120),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06892__B1 (.DIODE(net121),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06888__B1 (.DIODE(net121),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06896__B1 (.DIODE(net121),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout120_A (.DIODE(net121),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06874__B1 (.DIODE(net121),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06876__B1 (.DIODE(net121),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout119_A (.DIODE(net121),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout121_A (.DIODE(net122),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06872__B1 (.DIODE(net122),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06878__B1 (.DIODE(net122),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06880__B1 (.DIODE(net122),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout117_A (.DIODE(net122),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06860__B1 (.DIODE(net122),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout118_A (.DIODE(net122),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07406__B1 (.DIODE(net123),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07418__B1 (.DIODE(net123),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07001__B1 (.DIODE(net123),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06999__B1 (.DIODE(net123),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06997__B1 (.DIODE(net123),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06995__B1 (.DIODE(net123),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06993__B1 (.DIODE(net123),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06991__B1 (.DIODE(net123),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06989__B1 (.DIODE(net123),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06960__B1 (.DIODE(net123),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06997__A2_N (.DIODE(net125),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06995__A2_N (.DIODE(net125),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06993__A2_N (.DIODE(net125),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06991__A2_N (.DIODE(net125),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07408__A2_N (.DIODE(net125),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07418__A2_N (.DIODE(net125),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06989__A2_N (.DIODE(net125),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06987__A2_N (.DIODE(net125),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06960__A2_N (.DIODE(net125),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06814__B (.DIODE(net125),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07414__A2_N (.DIODE(net126),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07412__A2_N (.DIODE(net126),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07410__A2_N (.DIODE(net126),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06856__A2 (.DIODE(net126),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07406__A2_N (.DIODE(net126),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06815__B (.DIODE(net126),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06999__A2_N (.DIODE(net126),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07001__A2_N (.DIODE(net126),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07416__A2_N (.DIODE(net126),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout125_A (.DIODE(net126),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07404__A2 (.DIODE(net127),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06858__A2 (.DIODE(net127),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout126_A (.DIODE(net127),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06844__A2 (.DIODE(net127),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06850__A2 (.DIODE(net127),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06852__A2 (.DIODE(net127),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06848__A2 (.DIODE(net127),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06846__A2 (.DIODE(net127),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06842__A2 (.DIODE(net127),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06854__A2 (.DIODE(net127),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06874__A2 (.DIODE(net128),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06876__A2 (.DIODE(net128),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06870__A2 (.DIODE(net128),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06840__A2 (.DIODE(net128),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06836__A2 (.DIODE(net128),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06834__A2 (.DIODE(net128),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06832__A2 (.DIODE(net128),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06830__A2 (.DIODE(net128),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06816__A2 (.DIODE(net128),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06838__A2 (.DIODE(net128),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06906__A2 (.DIODE(net129),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06904__A2 (.DIODE(net129),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06894__A2 (.DIODE(net129),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06896__A2 (.DIODE(net129),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06900__A2 (.DIODE(net129),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06826__A2 (.DIODE(net129),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06822__A2 (.DIODE(net129),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06828__A2 (.DIODE(net129),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06824__A2 (.DIODE(net129),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06820__A2 (.DIODE(net129),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06880__A2 (.DIODE(net130),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06882__A2 (.DIODE(net130),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06884__A2 (.DIODE(net130),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06892__A2 (.DIODE(net130),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06890__A2 (.DIODE(net130),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06888__A2 (.DIODE(net130),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06902__A2 (.DIODE(net130),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06908__A2 (.DIODE(net130),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06898__A2 (.DIODE(net130),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout129_A (.DIODE(net130),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06886__A2 (.DIODE(net131),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout130_A (.DIODE(net131),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06818__A2 (.DIODE(net131),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06872__A2 (.DIODE(net131),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06878__A2 (.DIODE(net131),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout128_A (.DIODE(net131),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07419__A2 (.DIODE(net133),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07003__C (.DIODE(net133),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06962__A2 (.DIODE(net133),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06927__A2 (.DIODE(net133),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06926__A2 (.DIODE(net133),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06925__A2 (.DIODE(net133),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06924__A2 (.DIODE(net133),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06929__A2 (.DIODE(net133),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06928__A2 (.DIODE(net133),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06923__A2 (.DIODE(net133),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06946__A2 (.DIODE(net135),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06950__A2 (.DIODE(net135),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06949__A2 (.DIODE(net135),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06914__A2 (.DIODE(net135),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06953__A2 (.DIODE(net135),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06955__A2 (.DIODE(net135),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06956__A2 (.DIODE(net135),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06957__A2 (.DIODE(net135),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06954__A2 (.DIODE(net135),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06952__A2 (.DIODE(net135),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06922__A2 (.DIODE(net137),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06916__A2 (.DIODE(net137),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06915__A2 (.DIODE(net137),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06917__A2 (.DIODE(net137),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06918__A2 (.DIODE(net137),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06940__A2 (.DIODE(net137),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06912__A2 (.DIODE(net137),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06921__A2 (.DIODE(net137),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06920__A2 (.DIODE(net137),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06919__A2 (.DIODE(net137),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06934__A2 (.DIODE(net138),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06937__A2 (.DIODE(net138),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06938__A2 (.DIODE(net138),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06936__A2 (.DIODE(net138),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06941__A2 (.DIODE(net138),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06939__A2 (.DIODE(net138),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06942__A2 (.DIODE(net138),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout136_A (.DIODE(net138),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout135_A (.DIODE(net138),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout137_A (.DIODE(net138),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06935__A2 (.DIODE(net139),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06943__A2 (.DIODE(net139),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout138_A (.DIODE(net139),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout133_A (.DIODE(net139),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout134_A (.DIODE(net139),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout140_A (.DIODE(net142),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout141_A (.DIODE(net142),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06961__B1 (.DIODE(net142),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06911__A2 (.DIODE(net142),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07002__B (.DIODE(net142),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05953__B1 (.DIODE(net144),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05952__B1 (.DIODE(net144),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout143_A (.DIODE(net144),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05933__B1 (.DIODE(net144),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05930__B1 (.DIODE(net144),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05941__B1 (.DIODE(net145),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05938__B1 (.DIODE(net145),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05940__B1 (.DIODE(net145),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05939__B1 (.DIODE(net145),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05937__B1 (.DIODE(net145),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05932__B1 (.DIODE(net145),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05934__B1 (.DIODE(net145),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05931__B1 (.DIODE(net145),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05942__B1 (.DIODE(net145),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05943__B1 (.DIODE(net145),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05946__B1 (.DIODE(net146),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05948__B1 (.DIODE(net146),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05945__B1 (.DIODE(net146),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05947__B1 (.DIODE(net146),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05949__B1 (.DIODE(net146),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05944__B1 (.DIODE(net146),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05935__B1 (.DIODE(net146),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05936__B1 (.DIODE(net146),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout145_A (.DIODE(net146),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05769__B1 (.DIODE(net147),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05770__B1 (.DIODE(net147),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05771__B1 (.DIODE(net147),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05766__B1 (.DIODE(net147),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05763__B1 (.DIODE(net147),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05775__B1 (.DIODE(net147),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05772__B1 (.DIODE(net147),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05773__B1 (.DIODE(net147),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05774__B1 (.DIODE(net147),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05776__B1 (.DIODE(net147),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07417__S (.DIODE(net148),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07402__S (.DIODE(net148),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07413__S (.DIODE(net148),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07000__A2 (.DIODE(net148),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06998__A2 (.DIODE(net148),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06996__A2 (.DIODE(net148),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06994__A2 (.DIODE(net148),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06992__A2 (.DIODE(net148),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06990__A2 (.DIODE(net148),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06988__A2 (.DIODE(net148),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07420__A2 (.DIODE(net149),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07407__S (.DIODE(net149),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07415__S (.DIODE(net149),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout148_A (.DIODE(net149),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06709__A2 (.DIODE(net149),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06961__A3 (.DIODE(net149),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06958__A_N (.DIODE(net149),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06813__A2 (.DIODE(net149),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06710__A2 (.DIODE(net149),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06959__A2 (.DIODE(net149),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07400__A2 (.DIODE(net150),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06857__S (.DIODE(net150),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06855__S (.DIODE(net150),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07405__S (.DIODE(net150),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07411__S (.DIODE(net150),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07409__S (.DIODE(net150),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout149_A (.DIODE(net150),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout150_A (.DIODE(net151),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06843__S (.DIODE(net151),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06847__S (.DIODE(net151),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06851__S (.DIODE(net151),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06849__S (.DIODE(net151),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06845__S (.DIODE(net151),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06841__S (.DIODE(net151),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06853__S (.DIODE(net151),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06869__S (.DIODE(net152),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06877__S (.DIODE(net152),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06873__S (.DIODE(net152),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06817__S (.DIODE(net152),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06839__S (.DIODE(net152),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06835__S (.DIODE(net152),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06833__S (.DIODE(net152),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06831__S (.DIODE(net152),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06829__S (.DIODE(net152),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06837__S (.DIODE(net152),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06903__S (.DIODE(net153),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06901__S (.DIODE(net153),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06893__S (.DIODE(net153),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06895__S (.DIODE(net153),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06899__S (.DIODE(net153),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06825__S (.DIODE(net153),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06821__S (.DIODE(net153),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06827__S (.DIODE(net153),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06823__S (.DIODE(net153),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06819__S (.DIODE(net153),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06879__S (.DIODE(net154),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06881__S (.DIODE(net154),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06883__S (.DIODE(net154),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06891__S (.DIODE(net154),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06887__S (.DIODE(net154),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06889__S (.DIODE(net154),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06905__S (.DIODE(net154),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06907__S (.DIODE(net154),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06897__S (.DIODE(net154),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout153_A (.DIODE(net154),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06885__S (.DIODE(net155),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout154_A (.DIODE(net155),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06875__S (.DIODE(net155),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06871__S (.DIODE(net155),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout152_A (.DIODE(net155),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06859__S (.DIODE(net156),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06863__S (.DIODE(net156),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06867__S (.DIODE(net156),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06865__S (.DIODE(net156),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06861__S (.DIODE(net156),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout155_A (.DIODE(net156),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06138__B1 (.DIODE(net157),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06136__B1 (.DIODE(net157),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06135__B1 (.DIODE(net157),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06134__B1 (.DIODE(net157),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06132__B1 (.DIODE(net157),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06133__B1 (.DIODE(net157),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06155__C1 (.DIODE(net157),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06151__B1 (.DIODE(net157),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06137__B1 (.DIODE(net157),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06131__B1 (.DIODE(net157),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05940__A2 (.DIODE(net158),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05939__A2 (.DIODE(net158),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05943__A2 (.DIODE(net158),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05935__A2 (.DIODE(net158),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05932__A2 (.DIODE(net158),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05931__A2 (.DIODE(net158),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05934__A2 (.DIODE(net158),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05929__B (.DIODE(net158),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05936__A2 (.DIODE(net158),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05937__A2 (.DIODE(net158),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05941__A2 (.DIODE(net159),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05942__A2 (.DIODE(net159),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05938__A2 (.DIODE(net159),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout158_A (.DIODE(net159),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05933__A2 (.DIODE(net159),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05930__A2 (.DIODE(net159),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05946__A2 (.DIODE(net161),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05948__A2 (.DIODE(net161),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05947__A2 (.DIODE(net161),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05945__A2 (.DIODE(net161),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05944__A2 (.DIODE(net161),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05949__A2 (.DIODE(net161),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout160_A (.DIODE(net161),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05952__A2 (.DIODE(net161),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05953__A2 (.DIODE(net161),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05765__A2 (.DIODE(net162),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05769__A2 (.DIODE(net162),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05770__A2 (.DIODE(net162),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05771__A2 (.DIODE(net162),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05762__B (.DIODE(net162),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05776__A2 (.DIODE(net162),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05775__A2 (.DIODE(net162),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05772__A2 (.DIODE(net162),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05773__A2 (.DIODE(net162),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05774__A2 (.DIODE(net162),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05550__A2 (.DIODE(net166),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06140__A2 (.DIODE(net166),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06139__A2 (.DIODE(net166),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06138__A2 (.DIODE(net166),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06136__A2 (.DIODE(net166),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06135__A2 (.DIODE(net166),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06134__A2 (.DIODE(net166),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06133__A2 (.DIODE(net166),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06132__A2 (.DIODE(net166),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06123__B (.DIODE(net166),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05556__A2 (.DIODE(net167),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05544__A2 (.DIODE(net167),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout166_A (.DIODE(net167),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout165_A (.DIODE(net167),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout164_A (.DIODE(net167),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout168_A (.DIODE(net170),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05695__A2 (.DIODE(net170),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05568__A2 (.DIODE(net170),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05719__A2 (.DIODE(net170),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05713__A2 (.DIODE(net170),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05731__A2 (.DIODE(net170),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05725__A2 (.DIODE(net170),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05707__A2 (.DIODE(net170),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05701__A2 (.DIODE(net170),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05689__A2 (.DIODE(net170),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05640__A2 (.DIODE(net171),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05616__A2 (.DIODE(net171),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05586__A2 (.DIODE(net171),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05562__A2 (.DIODE(net171),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05646__A2 (.DIODE(net171),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout170_A (.DIODE(net171),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout169_A (.DIODE(net171),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08223__C1 (.DIODE(net172),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08349__C1 (.DIODE(net172),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08217__C1 (.DIODE(net172),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08221__C1 (.DIODE(net172),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08153__C1 (.DIODE(net172),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08152__A2 (.DIODE(net172),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08149__B (.DIODE(net172),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08145__A1 (.DIODE(net172),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08134__B1 (.DIODE(net172),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08128__C1 (.DIODE(net172),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout172_A (.DIODE(net174),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout173_A (.DIODE(net174),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08215__C1 (.DIODE(net174),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08157__C1 (.DIODE(net174),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08405__B1 (.DIODE(net174),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08283__C1 (.DIODE(net174),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08287__C1 (.DIODE(net174),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08155__C1 (.DIODE(net174),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08361__C1 (.DIODE(net176),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08363__C1 (.DIODE(net176),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08165__C1 (.DIODE(net176),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08357__C1 (.DIODE(net176),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08355__C1 (.DIODE(net176),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08167__C1 (.DIODE(net176),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08231__C1 (.DIODE(net176),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08229__C1 (.DIODE(net176),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08345__C1 (.DIODE(net176),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08353__C1 (.DIODE(net176),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08169__C1 (.DIODE(net177),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08365__C1 (.DIODE(net177),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08359__C1 (.DIODE(net177),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout176_A (.DIODE(net177),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08277__C1 (.DIODE(net177),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08341__C1 (.DIODE(net177),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08213__C1 (.DIODE(net177),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08293__C1 (.DIODE(net177),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout175_A (.DIODE(net177),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout185_A (.DIODE(net189),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout188_A (.DIODE(net189),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout179_A (.DIODE(net189),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout181_A (.DIODE(net189),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout180_A (.DIODE(net189),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08218__A2 (.DIODE(net190),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08228__A2 (.DIODE(net190),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08352__A2 (.DIODE(net190),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08226__A2 (.DIODE(net190),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08154__A2 (.DIODE(net190),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08151__B (.DIODE(net190),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08148__S (.DIODE(net190),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08138__B (.DIODE(net190),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08136__B1 (.DIODE(net190),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08224__A2 (.DIODE(net190),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout190_A (.DIODE(net192),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout191_A (.DIODE(net192),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08216__A2 (.DIODE(net192),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08288__A2 (.DIODE(net192),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08406__A2 (.DIODE(net192),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08156__A2 (.DIODE(net192),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08158__A2 (.DIODE(net192),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08284__A2 (.DIODE(net192),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08366__A2 (.DIODE(net194),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08166__A2 (.DIODE(net194),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08356__A2 (.DIODE(net194),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08168__A2 (.DIODE(net194),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08358__A2 (.DIODE(net194),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08354__A2 (.DIODE(net194),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08232__A2 (.DIODE(net194),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08230__A2 (.DIODE(net194),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08346__A2 (.DIODE(net194),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08350__A2 (.DIODE(net194),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08364__A2 (.DIODE(net195),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08170__A2 (.DIODE(net195),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08362__A2 (.DIODE(net195),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08360__A2 (.DIODE(net195),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout194_A (.DIODE(net195),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08296__A2 (.DIODE(net195),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08278__A2 (.DIODE(net195),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08342__A2 (.DIODE(net195),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08214__A2 (.DIODE(net195),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout193_A (.DIODE(net195),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08394__A2 (.DIODE(net197),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout196_A (.DIODE(net197),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08398__A2 (.DIODE(net197),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08402__A2 (.DIODE(net197),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08304__A2 (.DIODE(net197),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08306__A2 (.DIODE(net197),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08404__A2 (.DIODE(net197),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08302__A2 (.DIODE(net197),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout203_A (.DIODE(net205),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout204_A (.DIODE(net205),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08378__A2 (.DIODE(net205),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08186__A2 (.DIODE(net205),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08250__A2 (.DIODE(net205),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08248__A2 (.DIODE(net205),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08376__A2 (.DIODE(net205),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout202_A (.DIODE(net206),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout205_A (.DIODE(net206),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout197_A (.DIODE(net206),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout199_A (.DIODE(net206),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout198_A (.DIODE(net206),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06150__C_N (.DIODE(net207),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06268__B2 (.DIODE(net207),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06186__B2 (.DIODE(net207),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06124__B1 (.DIODE(net207),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06122__B1 (.DIODE(net207),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05538__B1 (.DIODE(net207),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05536__A_N (.DIODE(net207),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06155__B2 (.DIODE(net207),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06244__B2 (.DIODE(net207),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06129__B2 (.DIODE(net207),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06313__B2 (.DIODE(net208),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06130__C (.DIODE(net208),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06377__B2 (.DIODE(net208),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06369__B2 (.DIODE(net208),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06354__B2 (.DIODE(net208),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06334__B2 (.DIODE(net208),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06293__B2 (.DIODE(net208),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06212__B2 (.DIODE(net208),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05586__B2 (.DIODE(net212),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout211_A (.DIODE(net212),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout210_A (.DIODE(net212),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout209_A (.DIODE(net212),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05707__B2 (.DIODE(net212),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout212_A (.DIODE(net213),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05562__B2 (.DIODE(net213),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05556__B2 (.DIODE(net213),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05550__B2 (.DIODE(net213),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05544__B2 (.DIODE(net213),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05535__B1 (.DIODE(net213),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09334__B1 (.DIODE(net214),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09341__B1 (.DIODE(net214),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09338__B1 (.DIODE(net214),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09339__B1 (.DIODE(net214),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09346__B1 (.DIODE(net214),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09344__B1 (.DIODE(net214),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09345__B1 (.DIODE(net214),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09343__B1 (.DIODE(net214),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09342__B1 (.DIODE(net214),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09335__B1 (.DIODE(net214),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09317__B1 (.DIODE(net215),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09316__B1 (.DIODE(net215),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09315__B1 (.DIODE(net215),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09347__B1 (.DIODE(net215),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09349__B1 (.DIODE(net215),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09351__B1 (.DIODE(net215),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09348__B1 (.DIODE(net215),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09352__B1 (.DIODE(net215),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09353__B1 (.DIODE(net215),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09350__B1 (.DIODE(net215),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09360__B1 (.DIODE(net218),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09327__B1 (.DIODE(net218),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09329__B1 (.DIODE(net218),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout217_A (.DIODE(net218),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09333__B1 (.DIODE(net218),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09332__B1 (.DIODE(net218),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09331__B1 (.DIODE(net218),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout216_A (.DIODE(net219),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout215_A (.DIODE(net219),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout218_A (.DIODE(net219),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09340__B1 (.DIODE(net219),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09337__B1 (.DIODE(net219),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09336__B1 (.DIODE(net219),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout214_A (.DIODE(net219),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09377__A2 (.DIODE(net221),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09338__A2 (.DIODE(net221),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09340__A2 (.DIODE(net221),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09336__A2 (.DIODE(net221),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09365__A2 (.DIODE(net221),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09403__A2 (.DIODE(net221),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09397__A2 (.DIODE(net221),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09391__A2 (.DIODE(net221),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09394__A2 (.DIODE(net221),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09388__A2 (.DIODE(net221),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout221_A (.DIODE(net223),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout222_A (.DIODE(net223),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09334__A2 (.DIODE(net223),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09339__A2 (.DIODE(net223),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09335__A2 (.DIODE(net223),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout220_A (.DIODE(net223),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09356__A2 (.DIODE(net225),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09357__A2 (.DIODE(net225),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout224_A (.DIODE(net225),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09347__A2 (.DIODE(net225),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09349__A2 (.DIODE(net225),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09351__A2 (.DIODE(net225),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09348__A2 (.DIODE(net225),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09352__A2 (.DIODE(net225),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09353__A2 (.DIODE(net225),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09350__A2 (.DIODE(net225),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09326__A2 (.DIODE(net226),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09328__A2 (.DIODE(net226),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09323__A2 (.DIODE(net226),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09330__A2 (.DIODE(net226),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09360__A2 (.DIODE(net226),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09327__A2 (.DIODE(net226),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09359__A2 (.DIODE(net226),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09331__A2 (.DIODE(net226),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09332__A2 (.DIODE(net226),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09333__A2 (.DIODE(net226),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09358__A2 (.DIODE(net227),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09355__A2 (.DIODE(net227),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09329__A2 (.DIODE(net227),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout226_A (.DIODE(net227),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09354__A2 (.DIODE(net227),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout225_A (.DIODE(net227),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09362__S (.DIODE(net228),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09379__B1 (.DIODE(net228),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09376__B1 (.DIODE(net228),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09390__B1 (.DIODE(net228),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09382__S (.DIODE(net228),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09370__B1 (.DIODE(net228),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09387__B1 (.DIODE(net228),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09385__A2 (.DIODE(net228),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09396__B1 (.DIODE(net228),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09399__B1 (.DIODE(net228),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09393__B1 (.DIODE(net229),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09373__B1 (.DIODE(net229),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09367__B1 (.DIODE(net229),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout228_A (.DIODE(net229),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09364__B1 (.DIODE(net229),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09402__B1 (.DIODE(net229),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09410__A2 (.DIODE(net229),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09407__S (.DIODE(net229),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09405__S (.DIODE(net229),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08503__S (.DIODE(net233),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout232_A (.DIODE(net233),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08464__S (.DIODE(net233),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout231_A (.DIODE(net233),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout230_A (.DIODE(net233),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08532__S (.DIODE(net234),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08470__S (.DIODE(net234),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08469__S (.DIODE(net234),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08531__S (.DIODE(net234),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08529__S (.DIODE(net234),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08530__S (.DIODE(net234),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08436__S (.DIODE(net234),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08437__S (.DIODE(net234),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08438__S (.DIODE(net234),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08534__S (.DIODE(net234),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08535__S (.DIODE(net235),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08537__S (.DIODE(net235),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08538__S (.DIODE(net235),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08474__S (.DIODE(net235),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08473__S (.DIODE(net235),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08439__S (.DIODE(net235),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08440__S (.DIODE(net235),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08442__S (.DIODE(net235),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08441__S (.DIODE(net235),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08539__S (.DIODE(net235),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08471__S (.DIODE(net236),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08472__S (.DIODE(net236),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08536__S (.DIODE(net236),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout235_A (.DIODE(net236),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08533__S (.DIODE(net236),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08467__S (.DIODE(net236),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08468__S (.DIODE(net236),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout234_A (.DIODE(net236),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08453__S (.DIODE(net241),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08485__S (.DIODE(net241),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08517__S (.DIODE(net241),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout240_A (.DIODE(net241),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout238_A (.DIODE(net241),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout244_A (.DIODE(net246),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout245_A (.DIODE(net246),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08478__S (.DIODE(net246),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08540__S (.DIODE(net246),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08477__S (.DIODE(net246),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08541__S (.DIODE(net246),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout243_A (.DIODE(net246),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout246_A (.DIODE(net247),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout241_A (.DIODE(net247),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout236_A (.DIODE(net247),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07874__B1 (.DIODE(net248),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07889__B1 (.DIODE(net248),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07884__B1 (.DIODE(net248),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07879__B1 (.DIODE(net248),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07854__B1 (.DIODE(net248),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07849__B1 (.DIODE(net248),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09183__A (.DIODE(net248),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07834__B1 (.DIODE(net248),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07844__B1 (.DIODE(net248),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07839__B1 (.DIODE(net248),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07954__B1 (.DIODE(net249),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07964__B1 (.DIODE(net249),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07969__B1 (.DIODE(net249),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07794__B1 (.DIODE(net249),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07809__B1 (.DIODE(net249),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07819__B1 (.DIODE(net249),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07814__B1 (.DIODE(net249),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07824__B1 (.DIODE(net249),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07829__B1 (.DIODE(net249),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07804__B1 (.DIODE(net249),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07914__B1 (.DIODE(net251),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07949__B1 (.DIODE(net251),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07789__B1 (.DIODE(net251),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07919__B1 (.DIODE(net251),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07934__B1 (.DIODE(net251),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07924__B1 (.DIODE(net251),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07784__B1 (.DIODE(net251),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07779__B1 (.DIODE(net251),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07944__B1 (.DIODE(net251),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07939__B1 (.DIODE(net251),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07929__B1 (.DIODE(net252),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07774__B1 (.DIODE(net252),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout251_A (.DIODE(net252),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07894__B1 (.DIODE(net252),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07799__B1 (.DIODE(net252),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07909__B1 (.DIODE(net252),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07769__B1 (.DIODE(net252),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07764__B1 (.DIODE(net252),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07899__B1 (.DIODE(net252),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07904__B1 (.DIODE(net252),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout250_A (.DIODE(net253),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout249_A (.DIODE(net253),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout252_A (.DIODE(net253),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07859__B1 (.DIODE(net253),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07864__B1 (.DIODE(net253),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07869__B1 (.DIODE(net253),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout248_A (.DIODE(net253),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07943__C1 (.DIODE(net260),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07828__C1 (.DIODE(net260),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07818__C1 (.DIODE(net260),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07823__C1 (.DIODE(net260),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07813__C1 (.DIODE(net260),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07808__C1 (.DIODE(net260),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07798__C1 (.DIODE(net260),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07803__C1 (.DIODE(net260),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07793__C1 (.DIODE(net260),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07888__C1 (.DIODE(net260),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07928__C1 (.DIODE(net263),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout262_A (.DIODE(net263),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07878__C1 (.DIODE(net263),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07893__C1 (.DIODE(net263),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07883__C1 (.DIODE(net263),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07898__C1 (.DIODE(net263),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07903__C1 (.DIODE(net263),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07762__C1 (.DIODE(net263),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07908__C1 (.DIODE(net263),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07871__S (.DIODE(net264),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07861__S (.DIODE(net264),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07881__S (.DIODE(net264),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07684__A2 (.DIODE(net264),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07708__A2 (.DIODE(net264),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07702__A2 (.DIODE(net264),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07696__A2 (.DIODE(net264),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07690__A2 (.DIODE(net264),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07678__A2 (.DIODE(net264),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07756__S (.DIODE(net264),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07876__S (.DIODE(net265),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout264_A (.DIODE(net265),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07851__S (.DIODE(net265),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07712__B1 (.DIODE(net265),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07660__B1 (.DIODE(net265),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07856__S (.DIODE(net265),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07831__S (.DIODE(net265),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09383__B1 (.DIODE(net265),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07961__S (.DIODE(net266),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07956__S (.DIODE(net266),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07936__S (.DIODE(net266),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07941__S (.DIODE(net266),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07951__S (.DIODE(net266),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07776__S (.DIODE(net266),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07791__S (.DIODE(net266),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07796__S (.DIODE(net266),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07821__S (.DIODE(net266),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07801__S (.DIODE(net266),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07931__S (.DIODE(net267),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07896__S (.DIODE(net267),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07946__S (.DIODE(net267),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07760__S (.DIODE(net267),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07921__S (.DIODE(net267),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07786__S (.DIODE(net267),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07916__S (.DIODE(net267),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07906__S (.DIODE(net267),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07981__S (.DIODE(net267),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout266_A (.DIODE(net267),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07344__A1 (.DIODE(net268),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07330__A1 (.DIODE(net268),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07320__A1 (.DIODE(net268),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07322__A1 (.DIODE(net268),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07314__A1 (.DIODE(net268),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07310__A1 (.DIODE(net268),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07308__A1 (.DIODE(net268),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07304__B1 (.DIODE(net268),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07302__A1 (.DIODE(net268),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07316__B1 (.DIODE(net268),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout268_A (.DIODE(net270),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout269_A (.DIODE(net270),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07275__A1 (.DIODE(net270),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07291__B1 (.DIODE(net270),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07289__A1 (.DIODE(net270),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07286__A1 (.DIODE(net270),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07284__A1 (.DIODE(net270),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07277__A1 (.DIODE(net270),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07270__B1 (.DIODE(net270),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07268__A1 (.DIODE(net270),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07386__A1 (.DIODE(net271),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07399__A2 (.DIODE(net271),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07391__A2 (.DIODE(net271),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07393__A2 (.DIODE(net271),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07395__A2 (.DIODE(net271),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07397__A2 (.DIODE(net271),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07254__A1 (.DIODE(net271),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07248__B1_N (.DIODE(net271),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07247__A3 (.DIODE(net271),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07260__A1 (.DIODE(net271),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07365__B1 (.DIODE(net272),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07360__B1 (.DIODE(net272),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07262__B1 (.DIODE(net272),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07256__B1 (.DIODE(net272),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07370__A1 (.DIODE(net272),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07372__B1 (.DIODE(net272),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07358__A1 (.DIODE(net272),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07384__B1 (.DIODE(net272),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07389__A1 (.DIODE(net272),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout271_A (.DIODE(net272),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07363__A1 (.DIODE(net273),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07378__B (.DIODE(net273),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07376__A1 (.DIODE(net273),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout272_A (.DIODE(net273),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout270_A (.DIODE(net273),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07346__A2 (.DIODE(net274),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07330__B1 (.DIODE(net274),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07320__B1 (.DIODE(net274),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07322__B1 (.DIODE(net274),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07314__B1 (.DIODE(net274),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07310__B1 (.DIODE(net274),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07308__B1 (.DIODE(net274),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07304__A2 (.DIODE(net274),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07302__B1 (.DIODE(net274),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07316__A2 (.DIODE(net274),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout274_A (.DIODE(net276),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout275_A (.DIODE(net276),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07275__B1 (.DIODE(net276),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07292__A2 (.DIODE(net276),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07286__B1 (.DIODE(net276),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07289__B1 (.DIODE(net276),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07284__B1 (.DIODE(net276),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07277__B1 (.DIODE(net276),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07271__A2 (.DIODE(net276),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07268__B1 (.DIODE(net276),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07384__A2 (.DIODE(net277),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07399__B1 (.DIODE(net277),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07397__B1 (.DIODE(net277),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07391__B1 (.DIODE(net277),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07393__B1 (.DIODE(net277),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07395__B1 (.DIODE(net277),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07254__B1 (.DIODE(net277),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07247__B1 (.DIODE(net277),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07249__B2 (.DIODE(net277),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07260__B1 (.DIODE(net277),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07360__A2 (.DIODE(net278),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07262__A2 (.DIODE(net278),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07256__A2 (.DIODE(net278),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07358__B1 (.DIODE(net278),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07372__A2 (.DIODE(net278),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07370__B1 (.DIODE(net278),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07379__A2 (.DIODE(net278),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07389__B1 (.DIODE(net278),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07386__B1 (.DIODE(net278),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout277_A (.DIODE(net278),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07365__A2 (.DIODE(net279),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07363__B1 (.DIODE(net279),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07376__B1 (.DIODE(net279),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout278_A (.DIODE(net279),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout276_A (.DIODE(net279),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07755__S (.DIODE(net281),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07870__S (.DIODE(net281),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07875__S (.DIODE(net281),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07860__S (.DIODE(net281),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07855__S (.DIODE(net281),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07880__S (.DIODE(net281),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07749__S (.DIODE(net281),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07701__S (.DIODE(net281),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout280_A (.DIODE(net281),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout281_A (.DIODE(net282),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07657__A2 (.DIODE(net282),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07850__S (.DIODE(net282),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07845__S (.DIODE(net282),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07830__S (.DIODE(net282),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07835__S (.DIODE(net282),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07840__S (.DIODE(net282),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07865__S (.DIODE(net282),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07666__C (.DIODE(net282),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07713__A2 (.DIODE(net282),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07935__S (.DIODE(net283),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07800__S (.DIODE(net283),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07790__S (.DIODE(net283),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07825__S (.DIODE(net283),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07815__S (.DIODE(net283),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07810__S (.DIODE(net283),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07820__S (.DIODE(net283),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07805__S (.DIODE(net283),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07795__S (.DIODE(net283),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07885__S (.DIODE(net283),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09182__A (.DIODE(net287),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07421__A (.DIODE(net287),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06814__A (.DIODE(net287),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08023__A (.DIODE(net287),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08017__C1 (.DIODE(net287),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07003__B (.DIODE(net287),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06966__B (.DIODE(net287),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06965__B (.DIODE(net287),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06963__B1 (.DIODE(net287),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06961__A2 (.DIODE(net287),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07533__S (.DIODE(net289),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07540__S (.DIODE(net289),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07518__S (.DIODE(net289),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07568__S (.DIODE(net289),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07553__S (.DIODE(net289),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07537__S (.DIODE(net289),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07522__S (.DIODE(net289),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07525__S (.DIODE(net289),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07571__S (.DIODE(net289),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07556__S (.DIODE(net289),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07564__S (.DIODE(net290),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07561__S (.DIODE(net290),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07546__S (.DIODE(net290),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07530__S (.DIODE(net290),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07515__S (.DIODE(net290),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07549__S (.DIODE(net290),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07570__S1 (.DIODE(net292),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07554__S1 (.DIODE(net292),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07535__S1 (.DIODE(net292),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07536__S1 (.DIODE(net292),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07551__S1 (.DIODE(net292),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07552__S1 (.DIODE(net292),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07567__S1 (.DIODE(net292),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07566__S1 (.DIODE(net292),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07520__S1 (.DIODE(net292),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07521__S1 (.DIODE(net292),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07514__S1 (.DIODE(net293),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07544__S1 (.DIODE(net293),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07559__S1 (.DIODE(net293),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07560__S1 (.DIODE(net293),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07531__S1 (.DIODE(net293),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07517__S1 (.DIODE(net293),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07532__S1 (.DIODE(net293),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07563__S1 (.DIODE(net293),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07562__S1 (.DIODE(net293),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07516__S1 (.DIODE(net293),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07528__S1 (.DIODE(net294),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07545__S1 (.DIODE(net294),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07513__S1 (.DIODE(net294),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout293_A (.DIODE(net294),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07555__S1 (.DIODE(net294),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07539__S1 (.DIODE(net294),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07538__S1 (.DIODE(net294),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07548__S1 (.DIODE(net294),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07547__S1 (.DIODE(net294),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07524__S1 (.DIODE(net294),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07529__S1 (.DIODE(net295),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout294_A (.DIODE(net295),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07523__S1 (.DIODE(net295),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07569__S1 (.DIODE(net295),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout292_A (.DIODE(net295),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06453__A1 (.DIODE(net298),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06450__A1 (.DIODE(net298),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06449__B (.DIODE(net298),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06444__B (.DIODE(net298),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06445__A1 (.DIODE(net298),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06452__B (.DIODE(net298),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06455__B (.DIODE(net298),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout297_A (.DIODE(net298),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06471__B1 (.DIODE(net298),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06469__A (.DIODE(net298),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06456__A1 (.DIODE(net299),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06461__A (.DIODE(net299),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06462__A2 (.DIODE(net299),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout298_A (.DIODE(net299),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06430__A2 (.DIODE(net299),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06432__S (.DIODE(net300),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06447__S (.DIODE(net300),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06438__S (.DIODE(net300),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06440__S (.DIODE(net300),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06467__S (.DIODE(net300),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06436__S (.DIODE(net300),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06485__B1 (.DIODE(net300),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06484__S (.DIODE(net300),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06464__S (.DIODE(net300),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06459__S (.DIODE(net300),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06429__C (.DIODE(net301),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06417__S (.DIODE(net301),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06414__A2 (.DIODE(net301),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06413__B1 (.DIODE(net301),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06411__S (.DIODE(net301),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06406__S (.DIODE(net301),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06419__S (.DIODE(net301),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06425__S (.DIODE(net301),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06422__S (.DIODE(net301),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06427__S (.DIODE(net301),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06010__A (.DIODE(net304),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08721__A (.DIODE(net304),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09135__C (.DIODE(net304),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout302_A (.DIODE(net304),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout303_A (.DIODE(net304),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05657__A2 (.DIODE(net307),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05651__B1 (.DIODE(net307),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05693__A2 (.DIODE(net307),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05724__A2 (.DIODE(net307),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05700__A2 (.DIODE(net307),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05688__A2 (.DIODE(net307),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05705__A2 (.DIODE(net307),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05711__A2 (.DIODE(net307),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05717__A2 (.DIODE(net307),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05670__A2 (.DIODE(net307),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05663__A2 (.DIODE(net308),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05675__A2 (.DIODE(net308),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05681__A2 (.DIODE(net308),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout307_A (.DIODE(net308),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05729__A2 (.DIODE(net308),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05564__B1 (.DIODE(net309),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05558__B1 (.DIODE(net309),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05727__B1 (.DIODE(net309),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05570__B1 (.DIODE(net309),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05552__B1 (.DIODE(net309),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05546__B1 (.DIODE(net309),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05540__B1 (.DIODE(net309),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05522__A2 (.DIODE(net309),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06304__B2 (.DIODE(net309),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06374__A2 (.DIODE(net309),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05667__B1 (.DIODE(net310),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05661__B1 (.DIODE(net310),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05648__B1 (.DIODE(net310),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05655__B1 (.DIODE(net310),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05630__B1 (.DIODE(net310),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05691__B1 (.DIODE(net310),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05697__B1 (.DIODE(net310),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05703__B1 (.DIODE(net310),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05685__B1 (.DIODE(net310),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05709__B1 (.DIODE(net310),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout310_A (.DIODE(net311),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05588__B1 (.DIODE(net311),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05624__B1 (.DIODE(net311),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05721__B1 (.DIODE(net311),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05715__B1 (.DIODE(net311),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05600__B1 (.DIODE(net311),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05618__B1 (.DIODE(net311),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05612__B1 (.DIODE(net311),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05606__B1 (.DIODE(net311),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05594__B1 (.DIODE(net311),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05642__B1 (.DIODE(net312),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05636__B1 (.DIODE(net312),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05673__B1 (.DIODE(net312),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05679__B1 (.DIODE(net312),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout311_A (.DIODE(net312),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05582__B1 (.DIODE(net312),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05576__B1 (.DIODE(net312),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout309_A (.DIODE(net312),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout316_A (.DIODE(net317),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout315_A (.DIODE(net317),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout314_A (.DIODE(net317),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout313_A (.DIODE(net317),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09148__C1 (.DIODE(net317),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08756__B1 (.DIODE(net323),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08746__B1 (.DIODE(net323),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08775__B1 (.DIODE(net323),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08742__B1 (.DIODE(net323),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09298__B1 (.DIODE(net323),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08763__A2 (.DIODE(net323),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08760__B1 (.DIODE(net323),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08766__B1 (.DIODE(net323),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09287__B1 (.DIODE(net323),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09292__B1 (.DIODE(net323),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08806__B1 (.DIODE(net324),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08736__B1 (.DIODE(net324),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08798__A2 (.DIODE(net324),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08739__A2 (.DIODE(net324),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08795__B1 (.DIODE(net324),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08783__B1 (.DIODE(net324),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08802__B1 (.DIODE(net324),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08790__B1 (.DIODE(net324),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08786__A2 (.DIODE(net324),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08732__B1 (.DIODE(net324),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08357__B1 (.DIODE(net330),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08359__B1 (.DIODE(net330),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08233__B1 (.DIODE(net330),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08173__B1 (.DIODE(net330),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08367__B1 (.DIODE(net330),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08365__B1 (.DIODE(net330),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08361__B1 (.DIODE(net330),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08363__B1 (.DIODE(net330),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08169__B1 (.DIODE(net330),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout329_A (.DIODE(net331),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout330_A (.DIODE(net331),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout327_A (.DIODE(net331),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08229__B1 (.DIODE(net331),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08167__B1 (.DIODE(net331),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout328_A (.DIODE(net331),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08243__B1 (.DIODE(net335),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08245__B1 (.DIODE(net335),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08181__B1 (.DIODE(net335),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08373__B1 (.DIODE(net335),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout334_A (.DIODE(net335),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout332_A (.DIODE(net335),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout333_A (.DIODE(net335),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout335_A (.DIODE(net341),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08259__B1 (.DIODE(net341),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout340_A (.DIODE(net341),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout338_A (.DIODE(net341),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout331_A (.DIODE(net341),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06001__S (.DIODE(net348),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05997__S (.DIODE(net348),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05990__S (.DIODE(net348),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout347_A (.DIODE(net348),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout346_A (.DIODE(net348),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05988__S (.DIODE(net348),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05989__S (.DIODE(net348),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05991__S (.DIODE(net348),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05880__S (.DIODE(net350),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05879__S (.DIODE(net350),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05878__S (.DIODE(net350),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05877__S (.DIODE(net350),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05875__S (.DIODE(net350),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05874__S (.DIODE(net350),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05873__S (.DIODE(net350),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05872__S (.DIODE(net350),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05871__S (.DIODE(net350),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05876__S (.DIODE(net350),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout350_A (.DIODE(net352),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout351_A (.DIODE(net352),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout349_A (.DIODE(net352),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05890__S (.DIODE(net352),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05889__S (.DIODE(net352),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout352_A (.DIODE(net353),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05870__S (.DIODE(net353),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05869__S (.DIODE(net353),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05868__S (.DIODE(net353),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05867__S (.DIODE(net353),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09116__A1 (.DIODE(net353),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05603__A2 (.DIODE(net354),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05609__A2 (.DIODE(net354),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05615__A2 (.DIODE(net354),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05566__A2 (.DIODE(net354),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05561__A2 (.DIODE(net354),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05590__B1 (.DIODE(net354),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05578__B1 (.DIODE(net354),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05573__A2 (.DIODE(net354),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05585__A2 (.DIODE(net354),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05596__B1 (.DIODE(net354),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout354_A (.DIODE(net356),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout355_A (.DIODE(net356),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09084__B1 (.DIODE(net356),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05650__B (.DIODE(net356),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05549__A2 (.DIODE(net356),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05528__A (.DIODE(net356),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05555__A2 (.DIODE(net356),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05543__A2 (.DIODE(net356),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05669__A2 (.DIODE(net357),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05730__A2 (.DIODE(net357),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05718__A2 (.DIODE(net357),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05712__A2 (.DIODE(net357),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05706__A2 (.DIODE(net357),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05699__A2 (.DIODE(net357),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05687__A2 (.DIODE(net357),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05676__A2 (.DIODE(net357),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05664__A2 (.DIODE(net357),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05723__A2 (.DIODE(net357),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05658__A2 (.DIODE(net358),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05644__A2 (.DIODE(net358),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05638__A2 (.DIODE(net358),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05682__A2 (.DIODE(net358),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05652__A2 (.DIODE(net358),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05632__A2 (.DIODE(net358),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05626__A2 (.DIODE(net358),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05620__A2 (.DIODE(net358),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05694__A2 (.DIODE(net358),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout357_A (.DIODE(net358),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout358_A (.DIODE(net359),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05602__A2 (.DIODE(net359),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05584__A2 (.DIODE(net359),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05578__A2 (.DIODE(net359),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05567__A2 (.DIODE(net359),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05572__A2 (.DIODE(net359),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05596__A2 (.DIODE(net359),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05590__A2 (.DIODE(net359),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05608__A2 (.DIODE(net359),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05614__A2 (.DIODE(net359),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout359_A (.DIODE(net360),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05560__A2 (.DIODE(net360),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05554__A2 (.DIODE(net360),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05548__A2 (.DIODE(net360),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05542__A2 (.DIODE(net360),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09129__A1 (.DIODE(net360),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09118__B1 (.DIODE(net360),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06378__C (.DIODE(net360),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05529__A3 (.DIODE(net360),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06320__A2 (.DIODE(net361),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06299__B1 (.DIODE(net361),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06164__A2 (.DIODE(net361),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06276__A2 (.DIODE(net361),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06130__B (.DIODE(net361),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05494__B2 (.DIODE(net361),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06208__A2 (.DIODE(net361),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09147__A2 (.DIODE(net361),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06222__A2 (.DIODE(net361),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06251__A2 (.DIODE(net361),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08996__S (.DIODE(net366),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout365_A (.DIODE(net366),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08998__S (.DIODE(net366),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09005__S (.DIODE(net366),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08993__S (.DIODE(net366),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08992__S (.DIODE(net366),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08991__S (.DIODE(net366),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08990__S (.DIODE(net366),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08989__S (.DIODE(net366),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout369_A (.DIODE(net370),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08221__A2 (.DIODE(net370),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08217__A2 (.DIODE(net370),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08215__A2 (.DIODE(net370),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08157__A2 (.DIODE(net370),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08405__A2 (.DIODE(net370),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08119__B (.DIODE(net370),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08155__A2 (.DIODE(net370),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08283__A2 (.DIODE(net370),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08363__A2 (.DIODE(net373),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08361__A2 (.DIODE(net373),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08167__A2 (.DIODE(net373),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08165__A2 (.DIODE(net373),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08355__A2 (.DIODE(net373),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08353__A2 (.DIODE(net373),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08231__A2 (.DIODE(net373),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08229__A2 (.DIODE(net373),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08345__A2 (.DIODE(net373),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08349__A2 (.DIODE(net373),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08169__A2 (.DIODE(net374),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08359__A2 (.DIODE(net374),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08357__A2 (.DIODE(net374),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout373_A (.DIODE(net374),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout371_A (.DIODE(net374),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout372_A (.DIODE(net374),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout380_A (.DIODE(net382),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout381_A (.DIODE(net382),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08315__A2 (.DIODE(net382),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08313__A2 (.DIODE(net382),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout379_A (.DIODE(net382),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout382_A (.DIODE(net386),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout385_A (.DIODE(net386),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout376_A (.DIODE(net386),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout378_A (.DIODE(net386),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout377_A (.DIODE(net386),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout389_A (.DIODE(net390),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07836__S (.DIODE(net390),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07841__S (.DIODE(net390),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07846__S (.DIODE(net390),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07866__S (.DIODE(net390),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09383__A2 (.DIODE(net390),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07660__A2 (.DIODE(net390),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07712__A2 (.DIODE(net390),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07911__S (.DIODE(net391),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07966__S (.DIODE(net391),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07971__S (.DIODE(net391),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07976__S (.DIODE(net391),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07986__S (.DIODE(net391),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07811__S (.DIODE(net391),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07806__S (.DIODE(net391),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07826__S (.DIODE(net391),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07816__S (.DIODE(net391),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07886__S (.DIODE(net391),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07926__S (.DIODE(net392),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07766__S (.DIODE(net392),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07901__S (.DIODE(net392),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07891__S (.DIODE(net392),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout391_A (.DIODE(net392),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout390_A (.DIODE(net392),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07569__S0 (.DIODE(net394),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07523__S0 (.DIODE(net394),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07554__S0 (.DIODE(net394),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07566__S0 (.DIODE(net394),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07567__S0 (.DIODE(net394),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07536__S0 (.DIODE(net394),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07535__S0 (.DIODE(net394),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06093__B (.DIODE(net394),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07520__S0 (.DIODE(net394),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07521__S0 (.DIODE(net394),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07544__S0 (.DIODE(net395),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07514__S0 (.DIODE(net395),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07559__S0 (.DIODE(net395),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07560__S0 (.DIODE(net395),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07563__S0 (.DIODE(net395),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07562__S0 (.DIODE(net395),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07516__S0 (.DIODE(net395),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07531__S0 (.DIODE(net395),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07517__S0 (.DIODE(net395),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07532__S0 (.DIODE(net395),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07545__S0 (.DIODE(net396),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07513__S0 (.DIODE(net396),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout395_A (.DIODE(net396),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07570__S0 (.DIODE(net396),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07539__S0 (.DIODE(net396),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07538__S0 (.DIODE(net396),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07555__S0 (.DIODE(net396),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07547__S0 (.DIODE(net396),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07548__S0 (.DIODE(net396),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07524__S0 (.DIODE(net396),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07528__S0 (.DIODE(net397),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07529__S0 (.DIODE(net397),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout396_A (.DIODE(net397),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07552__S0 (.DIODE(net397),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07551__S0 (.DIODE(net397),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout394_A (.DIODE(net397),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout400_A (.DIODE(net401),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09402__A2 (.DIODE(net401),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09401__A (.DIODE(net401),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09406__S (.DIODE(net401),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09404__S (.DIODE(net401),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09364__A2 (.DIODE(net401),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09363__A (.DIODE(net401),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09383__C1 (.DIODE(net401),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05830__C (.DIODE(net401),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08775__A2 (.DIODE(net402),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05782__D (.DIODE(net402),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08861__A1 (.DIODE(net402),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05781__B (.DIODE(net402),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08760__A2 (.DIODE(net402),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08764__A2 (.DIODE(net402),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08766__A2 (.DIODE(net402),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09292__A2 (.DIODE(net402),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09287__A2 (.DIODE(net402),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08864__B (.DIODE(net402),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08825__A2 (.DIODE(net404),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08806__A2 (.DIODE(net404),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08799__A2 (.DIODE(net404),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08736__A2 (.DIODE(net404),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08795__A2 (.DIODE(net404),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08802__A2 (.DIODE(net404),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08790__A2 (.DIODE(net404),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08785__B (.DIODE(net404),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08783__A2 (.DIODE(net404),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08732__A2 (.DIODE(net404),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08740__A2 (.DIODE(net405),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08754__A2 (.DIODE(net405),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08810__A2 (.DIODE(net405),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08821__A2 (.DIODE(net405),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08817__A2 (.DIODE(net405),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08814__A2 (.DIODE(net405),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06356__A1 (.DIODE(net406),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06318__A2 (.DIODE(net406),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06248__A2 (.DIODE(net406),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06317__A (.DIODE(net406),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06958__C (.DIODE(net406),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06126__B1 (.DIODE(net406),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08019__A2 (.DIODE(net406),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08016__A (.DIODE(net406),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05744__B1 (.DIODE(net406),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09154__B2 (.DIODE(net406),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06153__A3 (.DIODE(net407),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07003__A (.DIODE(net407),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06130__D (.DIODE(net407),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06961__A1 (.DIODE(net407),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06370__A3 (.DIODE(net407),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06338__A1 (.DIODE(net407),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05730__B1 (.DIODE(net408),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05718__B1 (.DIODE(net408),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05712__B1 (.DIODE(net408),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05706__B1 (.DIODE(net408),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05694__B1 (.DIODE(net408),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05687__B1 (.DIODE(net408),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05669__B1 (.DIODE(net408),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05676__B1 (.DIODE(net408),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05664__B1 (.DIODE(net408),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05723__B1 (.DIODE(net408),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05658__B1 (.DIODE(net409),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05652__B1 (.DIODE(net409),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05682__B1 (.DIODE(net409),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05633__A2 (.DIODE(net409),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05627__A2 (.DIODE(net409),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05638__B1 (.DIODE(net409),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05644__B1 (.DIODE(net409),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05699__B1 (.DIODE(net409),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout408_A (.DIODE(net409),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05620__B1 (.DIODE(net410),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05591__A2 (.DIODE(net410),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05584__B1 (.DIODE(net410),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05608__B1 (.DIODE(net410),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05602__B1 (.DIODE(net410),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05573__B1 (.DIODE(net410),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05579__A2 (.DIODE(net410),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05597__A2 (.DIODE(net410),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05614__B1 (.DIODE(net410),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05566__B1 (.DIODE(net410),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout409_A (.DIODE(net411),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout410_A (.DIODE(net411),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05528__B (.DIODE(net411),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05865__B1 (.DIODE(net411),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05560__B1 (.DIODE(net411),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05554__B1 (.DIODE(net411),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05548__B1 (.DIODE(net411),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05542__B1 (.DIODE(net411),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05475__A2 (.DIODE(net414),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05486__A2 (.DIODE(net414),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05482__A2 (.DIODE(net414),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout413_A (.DIODE(net414),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05464__A2 (.DIODE(net414),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05461__A2 (.DIODE(net414),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05459__A2 (.DIODE(net414),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05455__A2 (.DIODE(net414),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05453__C (.DIODE(net414),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05463__A2 (.DIODE(net414),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07878__A1 (.DIODE(net417),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07873__A1 (.DIODE(net417),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07863__A1 (.DIODE(net417),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05816__B (.DIODE(net417),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07848__A1 (.DIODE(net417),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07713__B1 (.DIODE(net417),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07843__A1 (.DIODE(net417),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07838__A1 (.DIODE(net417),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07833__A1 (.DIODE(net417),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07853__A1 (.DIODE(net417),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07958__A1 (.DIODE(net418),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07953__A1 (.DIODE(net418),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07938__A1 (.DIODE(net418),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07803__A1 (.DIODE(net418),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07793__A1 (.DIODE(net418),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07818__A1 (.DIODE(net418),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07828__A1 (.DIODE(net418),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07813__A1 (.DIODE(net418),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07808__A1 (.DIODE(net418),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07823__A1 (.DIODE(net418),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout419_A (.DIODE(net422),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout418_A (.DIODE(net422),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout421_A (.DIODE(net422),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07773__A1 (.DIODE(net422),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07858__A1 (.DIODE(net422),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07868__A1 (.DIODE(net422),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08904__B (.DIODE(net422),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout417_A (.DIODE(net422),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08037__B1 (.DIODE(net423),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07607__B1 (.DIODE(net423),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07606__B (.DIODE(net423),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06096__B (.DIODE(net423),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09306__B1 (.DIODE(net423),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08845__B1 (.DIODE(net423),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08842__A1 (.DIODE(net423),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05778__A (.DIODE(net423),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05777__A (.DIODE(net423),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09092__A2 (.DIODE(net423),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08743__A1 (.DIODE(net425),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08749__A (.DIODE(net425),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08759__A (.DIODE(net425),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08751__A (.DIODE(net425),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08728__A (.DIODE(net425),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09296__A (.DIODE(net425),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08767__A1 (.DIODE(net425),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09286__A (.DIODE(net425),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09291__A (.DIODE(net425),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08763__B2 (.DIODE(net425),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08813__A (.DIODE(net426),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08809__B2 (.DIODE(net426),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08798__B2 (.DIODE(net426),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08796__A1 (.DIODE(net426),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08735__A (.DIODE(net426),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08782__A (.DIODE(net426),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08801__A (.DIODE(net426),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08791__A1 (.DIODE(net426),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08786__B2 (.DIODE(net426),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08731__A (.DIODE(net426),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout426_A (.DIODE(net428),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout427_A (.DIODE(net428),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08745__A (.DIODE(net428),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08757__A1 (.DIODE(net428),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout425_A (.DIODE(net428),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08786__C1 (.DIODE(net429),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08790__C1 (.DIODE(net429),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08736__C1 (.DIODE(net429),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08742__C1 (.DIODE(net429),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08766__C1 (.DIODE(net429),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09298__C1 (.DIODE(net429),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09292__C1 (.DIODE(net429),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09287__C1 (.DIODE(net429),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08769__B2 (.DIODE(net429),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08771__B2 (.DIODE(net429),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08824__C1 (.DIODE(net430),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08733__A1 (.DIODE(net430),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08817__C1 (.DIODE(net430),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08809__C1 (.DIODE(net430),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08814__C1 (.DIODE(net430),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08774__A (.DIODE(net430),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08831__A1 (.DIODE(net430),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07834__A1 (.DIODE(net431),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07839__A1 (.DIODE(net431),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07667__B2 (.DIODE(net431),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07869__A1 (.DIODE(net431),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07993__A1 (.DIODE(net431),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06593__A (.DIODE(net431),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05818__B (.DIODE(net431),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05817__B (.DIODE(net431),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07763__A (.DIODE(net431),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08719__A1 (.DIODE(net431),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07711__B2 (.DIODE(net432),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07699__B2 (.DIODE(net432),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07724__B2 (.DIODE(net432),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07705__B2 (.DIODE(net432),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07742__B2 (.DIODE(net432),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07736__B2 (.DIODE(net432),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07693__B2 (.DIODE(net432),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07687__B2 (.DIODE(net432),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07864__A1 (.DIODE(net432),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07859__A1 (.DIODE(net432),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07758__A1 (.DIODE(net433),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout432_A (.DIODE(net433),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07730__B2 (.DIODE(net433),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07664__A (.DIODE(net433),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07748__B2 (.DIODE(net433),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07754__B2 (.DIODE(net433),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07681__B2 (.DIODE(net433),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout433_A (.DIODE(net434),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07854__A1 (.DIODE(net434),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07849__A1 (.DIODE(net434),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07844__A1 (.DIODE(net434),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout431_A (.DIODE(net434),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07944__A1 (.DIODE(net435),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07804__A1 (.DIODE(net435),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07824__A1 (.DIODE(net435),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07814__A1 (.DIODE(net435),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07809__A1 (.DIODE(net435),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07799__A1 (.DIODE(net435),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07829__A1 (.DIODE(net435),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07819__A1 (.DIODE(net435),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07794__A1 (.DIODE(net435),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07889__A1 (.DIODE(net435),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07924__A1 (.DIODE(net438),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout437_A (.DIODE(net438),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07904__A1 (.DIODE(net438),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07764__A1 (.DIODE(net438),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07894__A1 (.DIODE(net438),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07899__A1 (.DIODE(net438),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07874__A1 (.DIODE(net438),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07884__A1 (.DIODE(net438),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07879__A1 (.DIODE(net438),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07909__A1 (.DIODE(net438),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06002__A (.DIODE(net439),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09143__C1 (.DIODE(net439),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06378__A (.DIODE(net439),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09066__A1 (.DIODE(net439),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05860__A (.DIODE(net439),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05529__A1 (.DIODE(net439),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05493__A (.DIODE(net439),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09110__A (.DIODE(net439),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05866__A (.DIODE(net439),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05917__A (.DIODE(net439),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09154__A1 (.DIODE(net440),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05515__A (.DIODE(net440),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05842__B (.DIODE(net440),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout439_A (.DIODE(net440),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05453__A (.DIODE(net440),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05287__A (.DIODE(net441),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_output72_A (.DIODE(net441),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__11886__A (.DIODE(net441),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__11885__A (.DIODE(net441),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__11884__A (.DIODE(net441),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__11883__A (.DIODE(net441),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__11882__A (.DIODE(net441),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__11797__D (.DIODE(net441),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06006__A (.DIODE(net441),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05538__A1 (.DIODE(net441),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout443_A (.DIODE(net444),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09114__A1 (.DIODE(net444),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09065__A1 (.DIODE(net444),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09008__A (.DIODE(net444),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06379__B (.DIODE(net444),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06127__A (.DIODE(net444),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06041__A (.DIODE(net444),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05797__A (.DIODE(net444),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05751__A (.DIODE(net444),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05510__A (.DIODE(net444),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05302__A (.DIODE(net448),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07994__A1 (.DIODE(net448),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05865__A1 (.DIODE(net448),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05841__B1 (.DIODE(net448),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06592__A (.DIODE(net448),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09141__C1 (.DIODE(net448),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05844__A (.DIODE(net448),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05836__A (.DIODE(net448),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09145__A1 (.DIODE(net448),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05526__A (.DIODE(net448),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07657__A1 (.DIODE(net449),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07665__A (.DIODE(net449),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08988__A (.DIODE(net449),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07718__A1 (.DIODE(net449),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07675__A1 (.DIODE(net449),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07671__A1 (.DIODE(net449),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08911__A (.DIODE(net449),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07714__B2 (.DIODE(net449),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout448_A (.DIODE(net449),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout451_A (.DIODE(net452),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09075__A1 (.DIODE(net452),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09139__A2 (.DIODE(net452),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09091__D_N (.DIODE(net452),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06003__B (.DIODE(net452),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05969__A (.DIODE(net452),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05968__A (.DIODE(net452),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08848__A (.DIODE(net452),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08842__C1 (.DIODE(net452),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05778__B (.DIODE(net452),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06347__C1 (.DIODE(net454),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06332__C1 (.DIODE(net454),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06303__C1 (.DIODE(net454),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06292__A1 (.DIODE(net454),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06256__C1 (.DIODE(net454),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06228__C1 (.DIODE(net454),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06154__A1 (.DIODE(net454),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05300__A (.DIODE(net454),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05795__A2 (.DIODE(net454),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout453_A (.DIODE(net454),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05749__B1 (.DIODE(net457),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05758__B (.DIODE(net457),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout456_A (.DIODE(net457),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05514__A1 (.DIODE(net457),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09073__A1 (.DIODE(net457),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09147__A1 (.DIODE(net457),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout455_A (.DIODE(net457),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09081__A2 (.DIODE(net459),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06300__B1 (.DIODE(net459),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09085__A1 (.DIODE(net459),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06967__A2 (.DIODE(net459),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06164__A1 (.DIODE(net459),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06163__A (.DIODE(net459),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06361__B1 (.DIODE(net459),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06252__B1 (.DIODE(net459),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06372__A (.DIODE(net459),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout458_A (.DIODE(net459),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09099__A1 (.DIODE(net462),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09070__A1 (.DIODE(net462),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09143__A1 (.DIODE(net462),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09097__A2 (.DIODE(net462),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09152__A2 (.DIODE(net462),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout460_A (.DIODE(net462),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout461_A (.DIODE(net462),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05583__B1 (.DIODE(net465),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05565__B1 (.DIODE(net465),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05559__B1 (.DIODE(net465),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05553__B1 (.DIODE(net465),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05547__B1 (.DIODE(net465),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05541__B1 (.DIODE(net465),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08969__A (.DIODE(net465),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06306__C1 (.DIODE(net465),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout464_A (.DIODE(net465),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout463_A (.DIODE(net465),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05577__B1 (.DIODE(net466),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout465_A (.DIODE(net466),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout462_A (.DIODE(net466),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08840__C (.DIODE(net466),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09140__A2 (.DIODE(net466),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09075__B2 (.DIODE(net466),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05657__B2 (.DIODE(net467),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05651__A1 (.DIODE(net467),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05613__B1 (.DIODE(net467),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05601__B1 (.DIODE(net467),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05589__B1 (.DIODE(net467),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05572__B2 (.DIODE(net467),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05607__B1 (.DIODE(net467),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05595__B1 (.DIODE(net467),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05619__B1 (.DIODE(net467),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05722__B1 (.DIODE(net467),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05643__B1 (.DIODE(net468),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05637__B1 (.DIODE(net468),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05631__B1 (.DIODE(net468),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05625__B1 (.DIODE(net468),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05668__B1 (.DIODE(net468),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05686__B1 (.DIODE(net468),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05698__B1 (.DIODE(net468),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05681__B2 (.DIODE(net468),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout467_A (.DIODE(net469),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout468_A (.DIODE(net469),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05729__B2 (.DIODE(net469),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05705__B2 (.DIODE(net469),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05693__B2 (.DIODE(net469),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05675__B2 (.DIODE(net469),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05663__B2 (.DIODE(net469),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05711__B2 (.DIODE(net469),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05717__B2 (.DIODE(net469),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07757__S (.DIODE(net475),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07710__A (.DIODE(net475),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07709__A (.DIODE(net475),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07877__A (.DIODE(net475),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07872__A (.DIODE(net475),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07862__A (.DIODE(net475),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07857__A (.DIODE(net475),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout474_A (.DIODE(net475),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07942__A (.DIODE(net476),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07827__A (.DIODE(net476),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07817__A (.DIODE(net476),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07797__A (.DIODE(net476),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07812__A (.DIODE(net476),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07807__A (.DIODE(net476),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07822__A (.DIODE(net476),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07802__A (.DIODE(net476),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07792__A (.DIODE(net476),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07887__A (.DIODE(net476),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07927__A (.DIODE(net478),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07947__A (.DIODE(net478),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07922__A (.DIODE(net478),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07892__A (.DIODE(net478),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07882__A (.DIODE(net478),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07897__A (.DIODE(net478),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07902__A (.DIODE(net478),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07767__A (.DIODE(net478),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07761__A (.DIODE(net478),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07907__A (.DIODE(net478),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout477_A (.DIODE(net480),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout476_A (.DIODE(net480),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout479_A (.DIODE(net480),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout478_A (.DIODE(net480),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout471_A (.DIODE(net480),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout475_A (.DIODE(net480),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07405__A0 (.DIODE(net482),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07422__B2 (.DIODE(net482),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06971__A (.DIODE(net482),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07004__B2 (.DIODE(net482),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06248__A1 (.DIODE(net482),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06222__A1 (.DIODE(net482),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06219__A (.DIODE(net482),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05490__B (.DIODE(net482),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05385__A (.DIODE(net482),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06988__B2 (.DIODE(net482),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08564__A1 (.DIODE(net491),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09220__A1 (.DIODE(net491),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09217__B1 (.DIODE(net491),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09242__B1 (.DIODE(net491),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09210__A1 (.DIODE(net491),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout490_A (.DIODE(net491),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08576__S1 (.DIODE(net492),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08607__S1 (.DIODE(net492),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08608__S1 (.DIODE(net492),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08578__S1 (.DIODE(net492),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08598__S1 (.DIODE(net492),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08599__S1 (.DIODE(net492),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08662__A1 (.DIODE(net492),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08661__A (.DIODE(net492),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08624__S1 (.DIODE(net492),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08625__S1 (.DIODE(net492),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08583__S1 (.DIODE(net494),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08590__S1 (.DIODE(net494),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08632__S1 (.DIODE(net494),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08631__S1 (.DIODE(net494),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08636__S1 (.DIODE(net494),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08595__S1 (.DIODE(net494),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08635__S1 (.DIODE(net494),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08594__S1 (.DIODE(net494),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08586__S1 (.DIODE(net494),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08585__S1 (.DIODE(net494),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08592__S1 (.DIODE(net495),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08581__S1 (.DIODE(net495),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08615__S1 (.DIODE(net495),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08616__S1 (.DIODE(net495),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout494_A (.DIODE(net495),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08573__S1 (.DIODE(net495),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08574__S1 (.DIODE(net495),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08620__S1 (.DIODE(net495),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08619__S1 (.DIODE(net495),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08596__S (.DIODE(net497),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08633__A (.DIODE(net497),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08584__A1 (.DIODE(net497),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08593__A1 (.DIODE(net497),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08637__S (.DIODE(net497),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08587__S (.DIODE(net497),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08621__S (.DIODE(net497),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08570__D (.DIODE(net498),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08569__B (.DIODE(net498),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08608__S0 (.DIODE(net498),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08607__S0 (.DIODE(net498),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08576__S0 (.DIODE(net498),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08578__S0 (.DIODE(net498),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08599__S0 (.DIODE(net498),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08598__S0 (.DIODE(net498),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08624__S0 (.DIODE(net498),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08625__S0 (.DIODE(net498),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08583__S0 (.DIODE(net500),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08590__S0 (.DIODE(net500),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08632__S0 (.DIODE(net500),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08631__S0 (.DIODE(net500),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08636__S0 (.DIODE(net500),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08595__S0 (.DIODE(net500),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08635__S0 (.DIODE(net500),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08594__S0 (.DIODE(net500),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08586__S0 (.DIODE(net500),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08585__S0 (.DIODE(net500),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08592__S0 (.DIODE(net501),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08581__S0 (.DIODE(net501),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08615__S0 (.DIODE(net501),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08616__S0 (.DIODE(net501),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout500_A (.DIODE(net501),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08573__S0 (.DIODE(net501),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08574__S0 (.DIODE(net501),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08620__S0 (.DIODE(net501),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08619__S0 (.DIODE(net501),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08753__C1 (.DIODE(net502),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08769__C1 (.DIODE(net502),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08771__C1 (.DIODE(net502),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08775__C1 (.DIODE(net502),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09303__S (.DIODE(net502),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09294__S (.DIODE(net502),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08860__A1 (.DIODE(net502),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08859__A (.DIODE(net502),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08856__B (.DIODE(net502),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05782__B (.DIODE(net502),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08778__C1 (.DIODE(net503),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05430__A (.DIODE(net503),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08804__B2 (.DIODE(net503),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08792__B1 (.DIODE(net503),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08795__C1 (.DIODE(net503),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08829__A1 (.DIODE(net503),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08830__A1 (.DIODE(net503),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08826__C1 (.DIODE(net503),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05782__C (.DIODE(net504),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08777__C1 (.DIODE(net504),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08861__B1 (.DIODE(net504),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05431__A (.DIODE(net504),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09302__S (.DIODE(net504),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09299__A1 (.DIODE(net504),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09293__A1 (.DIODE(net504),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09288__A1 (.DIODE(net504),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08760__C1 (.DIODE(net504),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08763__C1 (.DIODE(net504),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08732__C1 (.DIODE(net505),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08819__A1 (.DIODE(net505),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08826__A1 (.DIODE(net505),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08821__C1 (.DIODE(net505),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08806__C1 (.DIODE(net505),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08778__B2 (.DIODE(net505),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08739__C1 (.DIODE(net505),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05781__A (.DIODE(net505),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08746__C1 (.DIODE(net505),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout504_A (.DIODE(net505),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08729__S1 (.DIODE(net506),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08747__S1 (.DIODE(net506),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05780__A (.DIODE(net506),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09301__S1 (.DIODE(net506),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09300__S1 (.DIODE(net506),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09297__S1 (.DIODE(net506),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09289__S1 (.DIODE(net506),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09284__S1 (.DIODE(net506),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08865__B1 (.DIODE(net506),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08761__S1 (.DIODE(net506),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08815__S1 (.DIODE(net507),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08811__S1 (.DIODE(net507),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08803__S1 (.DIODE(net507),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08788__S1 (.DIODE(net507),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08737__S1 (.DIODE(net507),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05432__A (.DIODE(net507),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08747__S0 (.DIODE(net508),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08758__S (.DIODE(net508),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08750__S (.DIODE(net508),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05780__B (.DIODE(net508),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09285__S (.DIODE(net508),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08729__S0 (.DIODE(net508),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08765__S (.DIODE(net508),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08761__S0 (.DIODE(net508),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08728__B (.DIODE(net508),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09284__S0 (.DIODE(net508),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08748__S (.DIODE(net509),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout508_A (.DIODE(net509),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08866__A1 (.DIODE(net509),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08863__A (.DIODE(net509),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09301__S0 (.DIODE(net509),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09300__S0 (.DIODE(net509),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09290__S (.DIODE(net509),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09289__S0 (.DIODE(net509),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09297__S0 (.DIODE(net509),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09295__S (.DIODE(net509),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08816__S (.DIODE(net510),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08812__S (.DIODE(net510),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08823__S (.DIODE(net510),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08797__S (.DIODE(net510),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08805__S (.DIODE(net510),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08781__S (.DIODE(net510),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08800__S (.DIODE(net510),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08788__S0 (.DIODE(net510),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08784__S (.DIODE(net510),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08789__S (.DIODE(net510),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08803__S0 (.DIODE(net511),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08737__S0 (.DIODE(net511),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08794__S (.DIODE(net511),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08730__S (.DIODE(net511),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08762__S (.DIODE(net511),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08808__S (.DIODE(net511),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08752__S (.DIODE(net511),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08815__S0 (.DIODE(net511),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08734__S (.DIODE(net511),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08738__S (.DIODE(net511),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout510_A (.DIODE(net512),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08820__S (.DIODE(net512),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08811__S0 (.DIODE(net512),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout511_A (.DIODE(net512),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08741__S (.DIODE(net512),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08755__S (.DIODE(net512),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08744__S (.DIODE(net512),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout509_A (.DIODE(net512),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09158__B (.DIODE(net516),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07579__A (.DIODE(net516),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout515_A (.DIODE(net516),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07646__B2 (.DIODE(net516),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07639__B2 (.DIODE(net516),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07632__B2 (.DIODE(net516),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07625__B2 (.DIODE(net516),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07619__B2 (.DIODE(net516),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07587__B2 (.DIODE(net516),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05426__A (.DIODE(net516),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07604__B (.DIODE(net521),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05909__A (.DIODE(net521),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07579__B (.DIODE(net521),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07652__A1 (.DIODE(net521),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07646__A1 (.DIODE(net521),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07639__A1 (.DIODE(net521),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07632__A1 (.DIODE(net521),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07625__A1 (.DIODE(net521),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07619__A1 (.DIODE(net521),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07587__A1 (.DIODE(net521),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05515__C (.DIODE(net527),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06128__B (.DIODE(net527),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05800__A2 (.DIODE(net527),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09096__B1 (.DIODE(net527),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09094__B1 (.DIODE(net527),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09088__A1 (.DIODE(net527),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05798__A3 (.DIODE(net527),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05797__B (.DIODE(net527),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05501__B (.DIODE(net527),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05502__B (.DIODE(net527),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05551__B1 (.DIODE(net528),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05546__A2 (.DIODE(net528),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05540__A2 (.DIODE(net528),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05727__A2 (.DIODE(net528),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05582__A2 (.DIODE(net528),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05558__A2 (.DIODE(net528),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout527_A (.DIODE(net528),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06374__A1 (.DIODE(net528),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05503__B (.DIODE(net528),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08988__B (.DIODE(net528),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05654__B1 (.DIODE(net529),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05661__A2 (.DIODE(net529),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05673__A2 (.DIODE(net529),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05666__B1 (.DIODE(net529),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05709__A2 (.DIODE(net529),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05703__A2 (.DIODE(net529),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05697__A2 (.DIODE(net529),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05691__A2 (.DIODE(net529),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05679__A2 (.DIODE(net529),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05685__A2 (.DIODE(net529),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout529_A (.DIODE(net530),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05624__A2 (.DIODE(net530),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05600__A2 (.DIODE(net530),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05618__A2 (.DIODE(net530),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05612__A2 (.DIODE(net530),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05606__A2 (.DIODE(net530),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05594__A2 (.DIODE(net530),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05715__A2 (.DIODE(net530),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05721__A2 (.DIODE(net530),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05588__A2 (.DIODE(net530),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05630__A2 (.DIODE(net531),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05648__A2 (.DIODE(net531),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05641__B1 (.DIODE(net531),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05636__A2 (.DIODE(net531),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout530_A (.DIODE(net531),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout531_A (.DIODE(net532),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05575__B1 (.DIODE(net532),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05570__A2 (.DIODE(net532),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05563__B1 (.DIODE(net532),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout528_A (.DIODE(net532),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05498__A1 (.DIODE(net535),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout534_A (.DIODE(net535),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06318__C1 (.DIODE(net535),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06358__C1 (.DIODE(net535),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05446__A (.DIODE(net535),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09155__B2 (.DIODE(net535),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout533_A (.DIODE(net535),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05760__B (.DIODE(net536),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05761__A2 (.DIODE(net536),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09153__B1 (.DIODE(net536),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05926__A (.DIODE(net536),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05526__B (.DIODE(net536),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05839__C (.DIODE(net536),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09093__B2 (.DIODE(net536),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05840__A2 (.DIODE(net536),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05969__B (.DIODE(net536),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05968__B (.DIODE(net536),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05575__A2 (.DIODE(net537),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05563__A2 (.DIODE(net537),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05569__B1 (.DIODE(net537),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05557__B1 (.DIODE(net537),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05551__A2 (.DIODE(net537),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09149__A1 (.DIODE(net537),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09086__B2 (.DIODE(net537),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05926__B (.DIODE(net537),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05503__A (.DIODE(net537),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05502__A (.DIODE(net537),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05581__B1 (.DIODE(net538),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05539__B1 (.DIODE(net538),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05545__B1 (.DIODE(net538),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05587__B1 (.DIODE(net538),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05726__B1 (.DIODE(net538),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05660__B1 (.DIODE(net539),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05708__B1 (.DIODE(net539),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05599__B1 (.DIODE(net539),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05617__B1 (.DIODE(net539),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05611__B1 (.DIODE(net539),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05605__B1 (.DIODE(net539),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05623__B1 (.DIODE(net539),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05593__B1 (.DIODE(net539),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05714__B1 (.DIODE(net539),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05720__B1 (.DIODE(net539),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05629__B1 (.DIODE(net540),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05684__B1 (.DIODE(net540),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05672__B1 (.DIODE(net540),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05678__B1 (.DIODE(net540),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05641__A2 (.DIODE(net540),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05635__B1 (.DIODE(net540),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05647__B1 (.DIODE(net540),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05654__A2 (.DIODE(net540),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05666__A2 (.DIODE(net540),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout539_A (.DIODE(net541),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout540_A (.DIODE(net541),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05702__B1 (.DIODE(net541),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05696__B1 (.DIODE(net541),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05690__B1 (.DIODE(net541),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05552__A2 (.DIODE(net546),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05569__A2 (.DIODE(net546),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05557__A2 (.DIODE(net546),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05545__A2 (.DIODE(net546),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05539__A2 (.DIODE(net546),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05726__A2 (.DIODE(net546),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05576__A2 (.DIODE(net546),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09098__A1 (.DIODE(net546),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09070__B2 (.DIODE(net546),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout545_A (.DIODE(net546),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05629__A2 (.DIODE(net547),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05642__A2 (.DIODE(net547),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05647__A2 (.DIODE(net547),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05623__A2 (.DIODE(net547),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05660__A2 (.DIODE(net547),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05655__A2 (.DIODE(net547),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05672__A2 (.DIODE(net547),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05667__A2 (.DIODE(net547),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05678__A2 (.DIODE(net547),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05684__A2 (.DIODE(net547),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout547_A (.DIODE(net548),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05587__A2 (.DIODE(net548),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05611__A2 (.DIODE(net548),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05605__A2 (.DIODE(net548),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05599__A2 (.DIODE(net548),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05714__A2 (.DIODE(net548),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05593__A2 (.DIODE(net548),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05617__A2 (.DIODE(net548),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05720__A2 (.DIODE(net548),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05708__A2 (.DIODE(net548),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05635__A2 (.DIODE(net549),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout548_A (.DIODE(net549),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05696__A2 (.DIODE(net549),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05702__A2 (.DIODE(net549),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05690__A2 (.DIODE(net549),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09549__B (.DIODE(net558),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09591__B (.DIODE(net558),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09592__B (.DIODE(net558),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10270__B (.DIODE(net558),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout557_A (.DIODE(net558),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10269__B (.DIODE(net558),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout556_A (.DIODE(net558),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09614__B (.DIODE(net561),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09594__B (.DIODE(net561),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09443__B (.DIODE(net561),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout560_A (.DIODE(net561),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout558_A (.DIODE(net561),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10459__B (.DIODE(net570),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10458__B (.DIODE(net570),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10142__B (.DIODE(net570),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09520__B (.DIODE(net570),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09516__B (.DIODE(net570),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09510__B (.DIODE(net570),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10391__B (.DIODE(net570),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout569_A (.DIODE(net570),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout567_A (.DIODE(net571),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10545__B (.DIODE(net571),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout564_A (.DIODE(net571),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout570_A (.DIODE(net571),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout554_A (.DIODE(net571),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout555_A (.DIODE(net571),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout553_A (.DIODE(net571),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout561_A (.DIODE(net571),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09574__B (.DIODE(net582),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09573__B (.DIODE(net582),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09527__B (.DIODE(net582),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09526__B (.DIODE(net582),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09427__B (.DIODE(net582),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09426__B (.DIODE(net582),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09424__B (.DIODE(net582),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10402__B (.DIODE(net582),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10403__B (.DIODE(net582),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout581_A (.DIODE(net582),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout583_A (.DIODE(net584),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout575_A (.DIODE(net584),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout577_A (.DIODE(net584),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09604__B (.DIODE(net584),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout576_A (.DIODE(net584),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10151__B (.DIODE(net588),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10153__B (.DIODE(net588),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10249__B (.DIODE(net588),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10493__B (.DIODE(net588),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout587_A (.DIODE(net588),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout585_A (.DIODE(net588),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout586_A (.DIODE(net588),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout609_A (.DIODE(net611),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10346__B (.DIODE(net611),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10345__B (.DIODE(net611),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout610_A (.DIODE(net611),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout608_A (.DIODE(net611),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout606_A (.DIODE(net612),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout611_A (.DIODE(net612),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout597_A (.DIODE(net612),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout594_A (.DIODE(net612),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout601_A (.DIODE(net612),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09771__B (.DIODE(net623),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09940__B (.DIODE(net623),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09941__B (.DIODE(net623),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout622_A (.DIODE(net623),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09675__B (.DIODE(net623),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09666__B (.DIODE(net623),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09570__B (.DIODE(net623),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09902__B (.DIODE(net628),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout627_A (.DIODE(net628),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09936__B (.DIODE(net628),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09907__B (.DIODE(net628),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09906__B (.DIODE(net628),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09904__B (.DIODE(net628),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09903__B (.DIODE(net628),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09800__B (.DIODE(net628),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09769__B (.DIODE(net628),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09768__B (.DIODE(net628),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout626_A (.DIODE(net629),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09935__B (.DIODE(net629),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout628_A (.DIODE(net629),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout623_A (.DIODE(net629),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout624_A (.DIODE(net629),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09947__B (.DIODE(net629),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09942__B (.DIODE(net629),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout621_A (.DIODE(net630),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout615_A (.DIODE(net630),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout616_A (.DIODE(net630),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout629_A (.DIODE(net630),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout612_A (.DIODE(net630),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout630_A (.DIODE(net631),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout571_A (.DIODE(net631),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout588_A (.DIODE(net631),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout592_A (.DIODE(net631),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout584_A (.DIODE(net631),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout640_A (.DIODE(net643),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout639_A (.DIODE(net643),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout642_A (.DIODE(net643),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout641_A (.DIODE(net643),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout638_A (.DIODE(net643),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout647_A (.DIODE(net651),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout650_A (.DIODE(net651),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout648_A (.DIODE(net651),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout649_A (.DIODE(net651),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout643_A (.DIODE(net651),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout660_A (.DIODE(net661),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout653_A (.DIODE(net661),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout652_A (.DIODE(net661),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout655_A (.DIODE(net661),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout654_A (.DIODE(net661),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10471__B (.DIODE(net665),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout664_A (.DIODE(net665),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10472__B (.DIODE(net665),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10098__B (.DIODE(net665),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10022__B (.DIODE(net665),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10021__B (.DIODE(net665),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10020__B (.DIODE(net665),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10016__B (.DIODE(net665),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10552__B (.DIODE(net667),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10089__B (.DIODE(net667),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09993__B (.DIODE(net667),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09992__B (.DIODE(net667),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10553__B (.DIODE(net667),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10551__B (.DIODE(net667),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10550__B (.DIODE(net667),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10547__B (.DIODE(net667),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09989__B (.DIODE(net667),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09983__B (.DIODE(net667),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10556__B (.DIODE(net669),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10555__B (.DIODE(net669),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout668_A (.DIODE(net669),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10091__B (.DIODE(net669),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10548__B (.DIODE(net669),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10549__B (.DIODE(net669),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout666_A (.DIODE(net669),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout665_A (.DIODE(net670),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout662_A (.DIODE(net670),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout663_A (.DIODE(net670),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout669_A (.DIODE(net670),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout661_A (.DIODE(net670),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout679_A (.DIODE(net680),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout672_A (.DIODE(net680),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout671_A (.DIODE(net680),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout674_A (.DIODE(net680),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout673_A (.DIODE(net680),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout686_A (.DIODE(net689),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout685_A (.DIODE(net689),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout688_A (.DIODE(net689),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09898__B (.DIODE(net689),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout682_A (.DIODE(net689),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout681_A (.DIODE(net689),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout684_A (.DIODE(net689),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout683_A (.DIODE(net689),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10562__B (.DIODE(net695),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10559__B (.DIODE(net695),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10558__B (.DIODE(net695),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09995__B (.DIODE(net695),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10572__B (.DIODE(net695),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10571__B (.DIODE(net695),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10569__B (.DIODE(net695),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10557__B (.DIODE(net695),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09994__B (.DIODE(net695),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09991__B (.DIODE(net695),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10563__B (.DIODE(net696),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10568__B (.DIODE(net696),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout695_A (.DIODE(net696),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10295__B (.DIODE(net696),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10293__B (.DIODE(net696),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09998__B (.DIODE(net696),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09997__B (.DIODE(net696),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09996__B (.DIODE(net696),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09684__B (.DIODE(net697),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10579__B (.DIODE(net697),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10567__B (.DIODE(net697),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10565__B (.DIODE(net697),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10564__B (.DIODE(net697),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10561__B (.DIODE(net697),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10560__B (.DIODE(net697),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10554__B (.DIODE(net697),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09780__B (.DIODE(net697),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09716__B (.DIODE(net697),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09852__B (.DIODE(net698),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09781__B (.DIODE(net698),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09749__B (.DIODE(net698),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09748__B (.DIODE(net698),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09717__B (.DIODE(net698),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09685__B (.DIODE(net698),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout696_A (.DIODE(net700),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout699_A (.DIODE(net700),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout697_A (.DIODE(net700),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout698_A (.DIODE(net700),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout694_A (.DIODE(net700),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09884__B (.DIODE(net702),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09859__B (.DIODE(net702),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09854__B (.DIODE(net702),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09853__B (.DIODE(net702),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09723__B (.DIODE(net702),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09861__B (.DIODE(net702),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout701_A (.DIODE(net702),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09751__B (.DIODE(net705),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09721__B (.DIODE(net705),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09720__B (.DIODE(net705),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09719__B (.DIODE(net705),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09885__B (.DIODE(net705),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09822__B (.DIODE(net705),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09821__B (.DIODE(net705),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09783__B (.DIODE(net705),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09687__B (.DIODE(net705),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09686__B (.DIODE(net705),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09889__B (.DIODE(net710),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09888__B (.DIODE(net710),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout709_A (.DIODE(net710),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout705_A (.DIODE(net710),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout707_A (.DIODE(net710),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout703_A (.DIODE(net711),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout704_A (.DIODE(net711),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout702_A (.DIODE(net711),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout710_A (.DIODE(net711),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout700_A (.DIODE(net711),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout689_A (.DIODE(net712),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout680_A (.DIODE(net712),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout711_A (.DIODE(net712),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout651_A (.DIODE(net712),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout670_A (.DIODE(net712),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05738__S (.DIODE(net715),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05737__S (.DIODE(net715),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05736__S (.DIODE(net715),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05735__S (.DIODE(net715),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05734__S (.DIODE(net715),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05733__S (.DIODE(net715),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05288__A (.DIODE(net715),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout714_A (.DIODE(net715),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09548__A (.DIODE(net722),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09547__A (.DIODE(net722),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10273__A (.DIODE(net722),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10272__A (.DIODE(net722),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10271__A (.DIODE(net722),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09543__A (.DIODE(net722),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09542__A (.DIODE(net722),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09541__A (.DIODE(net722),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09540__A (.DIODE(net722),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09539__A (.DIODE(net722),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09549__A (.DIODE(net723),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09591__A (.DIODE(net723),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09592__A (.DIODE(net723),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10270__A (.DIODE(net723),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout722_A (.DIODE(net723),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10269__A (.DIODE(net723),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout721_A (.DIODE(net723),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09614__A (.DIODE(net726),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09594__A (.DIODE(net726),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09443__A (.DIODE(net726),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout725_A (.DIODE(net726),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout723_A (.DIODE(net726),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10459__A (.DIODE(net735),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10458__A (.DIODE(net735),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10142__A (.DIODE(net735),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09520__A (.DIODE(net735),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09516__A (.DIODE(net735),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09510__A (.DIODE(net735),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10391__A (.DIODE(net735),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout734_A (.DIODE(net735),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout732_A (.DIODE(net736),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10545__A (.DIODE(net736),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout729_A (.DIODE(net736),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout735_A (.DIODE(net736),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout719_A (.DIODE(net736),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout720_A (.DIODE(net736),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout718_A (.DIODE(net736),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout726_A (.DIODE(net736),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10416__A (.DIODE(net737),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10414__A (.DIODE(net737),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09546__A (.DIODE(net737),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10594__A (.DIODE(net737),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10590__A (.DIODE(net737),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09551__A (.DIODE(net737),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09550__A (.DIODE(net737),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09545__A (.DIODE(net737),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09544__A (.DIODE(net737),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09538__A (.DIODE(net737),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout738_A (.DIODE(net740),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout739_A (.DIODE(net740),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10417__A (.DIODE(net740),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10418__A (.DIODE(net740),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10419__A (.DIODE(net740),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout737_A (.DIODE(net740),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09574__A (.DIODE(net747),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09573__A (.DIODE(net747),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09527__A (.DIODE(net747),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09526__A (.DIODE(net747),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09427__A (.DIODE(net747),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09426__A (.DIODE(net747),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09424__A (.DIODE(net747),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10402__A (.DIODE(net747),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10403__A (.DIODE(net747),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout746_A (.DIODE(net747),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10392__A (.DIODE(net748),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10393__A (.DIODE(net748),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout747_A (.DIODE(net748),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout744_A (.DIODE(net748),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout743_A (.DIODE(net748),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout745_A (.DIODE(net748),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09582__A (.DIODE(net748),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout748_A (.DIODE(net749),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout740_A (.DIODE(net749),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout742_A (.DIODE(net749),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09604__A (.DIODE(net749),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout741_A (.DIODE(net749),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10151__A (.DIODE(net753),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10153__A (.DIODE(net753),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10249__A (.DIODE(net753),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10493__A (.DIODE(net753),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout752_A (.DIODE(net753),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout750_A (.DIODE(net753),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout751_A (.DIODE(net753),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout764_A (.DIODE(net766),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout765_A (.DIODE(net766),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10425__A (.DIODE(net766),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10460__A (.DIODE(net766),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout763_A (.DIODE(net766),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout770_A (.DIODE(net771),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09953__A (.DIODE(net771),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09954__A (.DIODE(net771),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09955__A (.DIODE(net771),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10612__A (.DIODE(net771),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout768_A (.DIODE(net771),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout771_A (.DIODE(net777),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout776_A (.DIODE(net777),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout762_A (.DIODE(net777),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout759_A (.DIODE(net777),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout766_A (.DIODE(net777),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09902__A (.DIODE(net793),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout792_A (.DIODE(net793),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09936__A (.DIODE(net793),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09907__A (.DIODE(net793),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09906__A (.DIODE(net793),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09904__A (.DIODE(net793),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09903__A (.DIODE(net793),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09800__A (.DIODE(net793),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09769__A (.DIODE(net793),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09768__A (.DIODE(net793),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout791_A (.DIODE(net794),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09935__A (.DIODE(net794),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout793_A (.DIODE(net794),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout788_A (.DIODE(net794),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout789_A (.DIODE(net794),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09947__A (.DIODE(net794),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09942__A (.DIODE(net794),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout786_A (.DIODE(net795),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout780_A (.DIODE(net795),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout781_A (.DIODE(net795),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout794_A (.DIODE(net795),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout777_A (.DIODE(net795),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout795_A (.DIODE(net796),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout736_A (.DIODE(net796),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout753_A (.DIODE(net796),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout757_A (.DIODE(net796),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout749_A (.DIODE(net796),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10231__A (.DIODE(net803),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10233__A (.DIODE(net803),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10454__A (.DIODE(net803),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10457__A (.DIODE(net803),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout802_A (.DIODE(net803),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout798_A (.DIODE(net803),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout797_A (.DIODE(net803),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout800_A (.DIODE(net803),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout799_A (.DIODE(net803),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout805_A (.DIODE(net808),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout804_A (.DIODE(net808),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout807_A (.DIODE(net808),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout806_A (.DIODE(net808),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout803_A (.DIODE(net808),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout812_A (.DIODE(net816),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout815_A (.DIODE(net816),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout813_A (.DIODE(net816),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout814_A (.DIODE(net816),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout808_A (.DIODE(net816),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10471__A (.DIODE(net830),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout829_A (.DIODE(net830),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10472__A (.DIODE(net830),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10098__A (.DIODE(net830),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10022__A (.DIODE(net830),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10021__A (.DIODE(net830),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10020__A (.DIODE(net830),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10016__A (.DIODE(net830),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10552__A (.DIODE(net832),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10089__A (.DIODE(net832),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09993__A (.DIODE(net832),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09992__A (.DIODE(net832),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10553__A (.DIODE(net832),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10551__A (.DIODE(net832),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10550__A (.DIODE(net832),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10547__A (.DIODE(net832),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09989__A (.DIODE(net832),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09983__A (.DIODE(net832),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10556__A (.DIODE(net834),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10555__A (.DIODE(net834),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout833_A (.DIODE(net834),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10091__A (.DIODE(net834),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10548__A (.DIODE(net834),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10549__A (.DIODE(net834),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout831_A (.DIODE(net834),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout830_A (.DIODE(net835),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout827_A (.DIODE(net835),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout828_A (.DIODE(net835),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout834_A (.DIODE(net835),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout826_A (.DIODE(net835),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10303__A (.DIODE(net844),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10304__A (.DIODE(net844),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout843_A (.DIODE(net844),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout840_A (.DIODE(net844),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout841_A (.DIODE(net844),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout844_A (.DIODE(net845),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout837_A (.DIODE(net845),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout836_A (.DIODE(net845),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout839_A (.DIODE(net845),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout838_A (.DIODE(net845),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout851_A (.DIODE(net854),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout850_A (.DIODE(net854),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout853_A (.DIODE(net854),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09898__A (.DIODE(net854),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout847_A (.DIODE(net854),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout846_A (.DIODE(net854),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout849_A (.DIODE(net854),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout848_A (.DIODE(net854),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10562__A (.DIODE(net860),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10559__A (.DIODE(net860),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10558__A (.DIODE(net860),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09995__A (.DIODE(net860),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10572__A (.DIODE(net860),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10571__A (.DIODE(net860),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10569__A (.DIODE(net860),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10557__A (.DIODE(net860),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09994__A (.DIODE(net860),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09991__A (.DIODE(net860),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09684__A (.DIODE(net862),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10579__A (.DIODE(net862),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10567__A (.DIODE(net862),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10565__A (.DIODE(net862),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10564__A (.DIODE(net862),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10561__A (.DIODE(net862),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10560__A (.DIODE(net862),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10554__A (.DIODE(net862),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09780__A (.DIODE(net862),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09716__A (.DIODE(net862),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout861_A (.DIODE(net865),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout864_A (.DIODE(net865),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout862_A (.DIODE(net865),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout863_A (.DIODE(net865),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout859_A (.DIODE(net865),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09751__A (.DIODE(net870),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09721__A (.DIODE(net870),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09720__A (.DIODE(net870),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09719__A (.DIODE(net870),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09885__A (.DIODE(net870),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09822__A (.DIODE(net870),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09821__A (.DIODE(net870),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09783__A (.DIODE(net870),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09687__A (.DIODE(net870),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09686__A (.DIODE(net870),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09889__A (.DIODE(net875),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09888__A (.DIODE(net875),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout874_A (.DIODE(net875),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout870_A (.DIODE(net875),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout872_A (.DIODE(net875),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout868_A (.DIODE(net876),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout869_A (.DIODE(net876),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout867_A (.DIODE(net876),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout875_A (.DIODE(net876),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout865_A (.DIODE(net876),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout854_A (.DIODE(net877),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout845_A (.DIODE(net877),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout876_A (.DIODE(net877),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout816_A (.DIODE(net877),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout835_A (.DIODE(net877),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_A (.DIODE(clknet_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_A (.DIODE(clknet_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_A (.DIODE(clknet_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_A (.DIODE(clknet_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_A (.DIODE(clknet_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_A (.DIODE(clknet_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_A (.DIODE(clknet_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_A (.DIODE(clknet_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_A (.DIODE(clknet_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_A (.DIODE(clknet_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_A (.DIODE(clknet_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_A (.DIODE(clknet_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_A (.DIODE(clknet_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_A (.DIODE(clknet_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_A (.DIODE(clknet_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_A (.DIODE(clknet_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_120_clk_A (.DIODE(clknet_4_0_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_119_clk_A (.DIODE(clknet_4_0_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_118_clk_A (.DIODE(clknet_4_0_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_117_clk_A (.DIODE(clknet_4_0_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_116_clk_A (.DIODE(clknet_4_0_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_clk_A (.DIODE(clknet_4_0_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_clk_A (.DIODE(clknet_4_0_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_clk_A (.DIODE(clknet_4_0_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_clk_A (.DIODE(clknet_4_1_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_clk_A (.DIODE(clknet_4_1_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_clk_A (.DIODE(clknet_4_1_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_clk_A (.DIODE(clknet_4_1_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_clk_A (.DIODE(clknet_4_1_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_clk_A (.DIODE(clknet_4_1_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_clk_A (.DIODE(clknet_4_1_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_clk_A (.DIODE(clknet_4_1_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_115_clk_A (.DIODE(clknet_4_2_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_114_clk_A (.DIODE(clknet_4_2_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_113_clk_A (.DIODE(clknet_4_2_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_112_clk_A (.DIODE(clknet_4_2_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_111_clk_A (.DIODE(clknet_4_2_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_110_clk_A (.DIODE(clknet_4_2_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_109_clk_A (.DIODE(clknet_4_2_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_108_clk_A (.DIODE(clknet_4_2_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_107_clk_A (.DIODE(clknet_4_3_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_106_clk_A (.DIODE(clknet_4_3_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_105_clk_A (.DIODE(clknet_4_3_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_clk_A (.DIODE(clknet_4_3_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_clk_A (.DIODE(clknet_4_3_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_clk_A (.DIODE(clknet_4_3_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_clk_A (.DIODE(clknet_4_4_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_clk_A (.DIODE(clknet_4_4_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_clk_A (.DIODE(clknet_4_4_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_clk_A (.DIODE(clknet_4_4_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_clk_A (.DIODE(clknet_4_4_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_clk_A (.DIODE(clknet_4_4_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_clk_A (.DIODE(clknet_4_4_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_clk_A (.DIODE(clknet_4_4_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_32_clk_A (.DIODE(clknet_4_5_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_clk_A (.DIODE(clknet_4_5_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_clk_A (.DIODE(clknet_4_5_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_clk_A (.DIODE(clknet_4_5_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_clk_A (.DIODE(clknet_4_5_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_clk_A (.DIODE(clknet_4_5_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_clk_A (.DIODE(clknet_4_5_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_43_clk_A (.DIODE(clknet_4_6_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_42_clk_A (.DIODE(clknet_4_6_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_41_clk_A (.DIODE(clknet_4_6_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_40_clk_A (.DIODE(clknet_4_6_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_clk_A (.DIODE(clknet_4_6_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_clk_A (.DIODE(clknet_4_6_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_clk_A (.DIODE(clknet_4_6_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_clk_A (.DIODE(clknet_4_6_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_39_clk_A (.DIODE(clknet_4_7_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_38_clk_A (.DIODE(clknet_4_7_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_37_clk_A (.DIODE(clknet_4_7_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_36_clk_A (.DIODE(clknet_4_7_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_35_clk_A (.DIODE(clknet_4_7_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_34_clk_A (.DIODE(clknet_4_7_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_33_clk_A (.DIODE(clknet_4_7_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_101_clk_A (.DIODE(clknet_4_8_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_100_clk_A (.DIODE(clknet_4_8_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_99_clk_A (.DIODE(clknet_4_8_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_98_clk_A (.DIODE(clknet_4_8_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_97_clk_A (.DIODE(clknet_4_8_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_96_clk_A (.DIODE(clknet_4_8_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_95_clk_A (.DIODE(clknet_4_8_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_104_clk_A (.DIODE(clknet_4_9_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_103_clk_A (.DIODE(clknet_4_9_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_102_clk_A (.DIODE(clknet_4_9_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_78_clk_A (.DIODE(clknet_4_9_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_77_clk_A (.DIODE(clknet_4_9_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_76_clk_A (.DIODE(clknet_4_9_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_75_clk_A (.DIODE(clknet_4_9_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_94_clk_A (.DIODE(clknet_4_10_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_93_clk_A (.DIODE(clknet_4_10_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_92_clk_A (.DIODE(clknet_4_10_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_91_clk_A (.DIODE(clknet_4_10_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_90_clk_A (.DIODE(clknet_4_10_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_89_clk_A (.DIODE(clknet_4_10_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_88_clk_A (.DIODE(clknet_4_10_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_87_clk_A (.DIODE(clknet_4_10_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_86_clk_A (.DIODE(clknet_4_10_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_85_clk_A (.DIODE(clknet_4_11_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_84_clk_A (.DIODE(clknet_4_11_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_83_clk_A (.DIODE(clknet_4_11_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_82_clk_A (.DIODE(clknet_4_11_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_81_clk_A (.DIODE(clknet_4_11_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_80_clk_A (.DIODE(clknet_4_11_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_79_clk_A (.DIODE(clknet_4_11_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_74_clk_A (.DIODE(clknet_4_12_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_73_clk_A (.DIODE(clknet_4_12_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_72_clk_A (.DIODE(clknet_4_12_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_71_clk_A (.DIODE(clknet_4_12_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_47_clk_A (.DIODE(clknet_4_12_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_46_clk_A (.DIODE(clknet_4_12_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_45_clk_A (.DIODE(clknet_4_12_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_44_clk_A (.DIODE(clknet_4_12_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_55_clk_A (.DIODE(clknet_4_13_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_54_clk_A (.DIODE(clknet_4_13_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_53_clk_A (.DIODE(clknet_4_13_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_52_clk_A (.DIODE(clknet_4_13_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_51_clk_A (.DIODE(clknet_4_13_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_50_clk_A (.DIODE(clknet_4_13_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_49_clk_A (.DIODE(clknet_4_13_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_48_clk_A (.DIODE(clknet_4_13_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_70_clk_A (.DIODE(clknet_4_14_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_69_clk_A (.DIODE(clknet_4_14_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_68_clk_A (.DIODE(clknet_4_14_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_67_clk_A (.DIODE(clknet_4_14_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_66_clk_A (.DIODE(clknet_4_14_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_65_clk_A (.DIODE(clknet_4_14_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_64_clk_A (.DIODE(clknet_4_14_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_63_clk_A (.DIODE(clknet_4_14_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_62_clk_A (.DIODE(clknet_4_15_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_61_clk_A (.DIODE(clknet_4_15_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_60_clk_A (.DIODE(clknet_4_15_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_59_clk_A (.DIODE(clknet_4_15_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_58_clk_A (.DIODE(clknet_4_15_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_57_clk_A (.DIODE(clknet_4_15_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_56_clk_A (.DIODE(clknet_4_15_0_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07924__B2 (.DIODE(net1559),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07363__B2 (.DIODE(net1559),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(ACK_I),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(DAT_I[10]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(DAT_I[18]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(DAT_I[24]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(DAT_I[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_01191_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_02725_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_03182_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_04146_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(_04150_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(en),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(gpio_in[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(gpio_in[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(gpio_in[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(gpio_in[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(\top.WB.CPU_DAT_O[19] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(\top.WB.CPU_DAT_O[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(\top.WB.CPU_DAT_O[24] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(\top.WB.CPU_DAT_O[27] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(\top.WB.CPU_DAT_O[28] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(\top.cb_syn.end_cnt[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(net253),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(net295),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(net353),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(net411),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(DAT_I[17]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(_04249_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(\top.WB.CPU_DAT_O[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(\top.WB.CPU_DAT_O[28] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(\top.cb_syn.end_cnt[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(_02735_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(\top.WB.CPU_DAT_O[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(\top.WB.CPU_DAT_O[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(\top.WB.CPU_DAT_O[28] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(net212),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_175 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_376 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_419 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_447 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_503 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_520 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_526 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_572 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_587 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_597 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_0_606 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_614 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_0_617 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_621 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_0_627 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_635 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_641 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_0_645 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_678 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_688 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_706 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_0_718 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_726 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_0_729 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_46 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_70 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_200 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_439 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_456 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_1_609 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_613 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_668 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_671 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_715 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_727 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_1_729 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_123 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_244 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_309 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_436 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_506 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_510 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_535 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_564 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_620 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_643 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_649 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_699 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_703 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_711 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_723 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_728 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_98 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_286 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_317 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_400 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_460 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_481 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_540 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_589 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_617 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_671 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_703 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_19 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_134 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_179 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_185 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_228 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_340 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_365 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_395 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_405 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_447 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_544 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_616 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_645 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_688 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_699 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_84 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_194 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_232 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_252 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_337 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_349 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_494 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_514 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_548 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_601 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_646 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_671 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_10 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_38 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_70 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_205 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_275 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_376 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_689 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_90 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_144 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_307 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_381 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_471 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_489 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_534 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_568 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_587 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_617 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_646 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_670 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_675 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_713 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_129 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_153 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_210 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_315 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_396 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_481 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_515 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_579 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_8_585 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_593 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_8_620 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_8_641 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_645 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_670 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_681 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_691 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_732 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_7 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_25 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_158 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_361 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_370 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_373 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_424 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_460 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_511 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_523 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_569 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_575 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_597 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_614 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_617 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_648 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_705 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_727 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_99 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_348 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_378 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_456 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_465 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_477 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_497 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_510 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_523 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_10_536 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_546 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_10_565 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_573 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_599 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_612 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_618 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_621 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_643 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_676 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_45 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_126 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_474 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_488 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_502 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_512 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_530 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_539 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_566 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_580 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_11_595 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_622 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_651 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_664 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_688 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_45 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_134 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_166 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_177 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_315 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_324 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_331 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_343 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_385 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_488 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_502 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_508 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_518 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_545 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_556 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_568 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_12_580 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_12_627 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_635 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_642 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_645 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_649 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_660 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_719 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_723 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_66 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_143 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_352 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_462 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_478 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_490 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_502 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_517 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_523 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_527 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_531 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_535 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_547 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_564 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_568 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_593 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_604 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_608 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_671 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_722 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_367 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_406 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_470 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_477 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_14_485 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_493 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_505 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_509 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_530 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_537 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_556 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_568 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_14_580 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_14_589 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_597 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_609 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_623 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_642 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_645 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_682 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_74 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_130 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_152 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_188 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_359 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_462 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_474 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_479 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_497 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_505 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_511 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_515 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_527 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_542 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_568 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_15_588 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_592 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_620 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_671 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_678 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_732 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_10 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_97 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_203 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_455 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_462 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_474 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_489 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_495 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_510 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_514 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_538 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_16_558 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_16_564 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_572 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_580 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_16_589 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_16_597 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_677 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_682 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_686 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_732 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_70 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_94 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_135 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_203 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_240 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_249 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_270 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_325 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_466 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_476 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_17_491 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_512 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_535 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_541 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_565 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_592 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_598 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_650 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_675 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_685 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_23 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_72 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_309 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_367 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_447 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_466 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_470 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_477 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_18_490 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_540 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_643 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_677 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_690 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_712 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_16 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_39 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_47 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_324 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_395 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_414 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_451 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_471 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_19_495 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_503 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_507 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_516 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_528 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_547 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_554 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_561 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_606 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_619 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_641 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_649 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_671 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_686 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_60 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_91 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_112 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_125 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_156 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_235 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_245 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_292 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_460 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_533 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_591 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_671 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_676 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_699 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_718 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_724 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_10 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_18 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_50 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_92 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_118 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_162 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_330 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_393 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_525 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_584 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_611 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_634 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_698 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_705 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_727 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_732 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_17 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_40 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_50 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_75 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_143 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_206 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_231 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_261 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_302 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_324 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_345 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_363 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_450 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_459 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_497 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_509 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_540 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_561 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_640 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_643 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_728 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_66 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_304 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_370 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_376 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_492 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_497 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_503 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_507 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_576 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_626 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_689 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_727 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_729 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_732 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_93 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_177 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_327 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_391 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_414 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_455 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_601 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_658 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_667 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_66 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_162 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_186 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_306 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_359 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_382 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_395 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_422 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_464 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_499 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_549 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_644 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_663 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_677 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_686 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_705 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_45 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_59 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_249 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_309 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_367 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_405 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_461 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_465 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_472 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_500 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_531 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_533 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_683 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_726 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_42 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_94 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_147 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_186 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_209 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_286 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_330 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_463 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_477 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_492 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_511 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_531 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_559 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_584 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_588 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_650 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_673 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_686 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_707 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_63 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_280 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_301 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_315 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_351 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_419 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_432 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_475 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_490 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_502 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_518 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_531 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_553 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_578 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_625 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_649 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_688 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_693 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_699 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_701 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_7 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_34 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_78 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_109 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_218 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_341 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_348 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_409 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_413 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_429 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_29_464 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_500 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_29_568 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_623 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_668 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_704 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_145 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_186 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_334 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_378 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_30_409 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_415 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_419 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_421 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_431 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_443 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_448 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_458 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_475 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_30_477 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_30_487 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_30_495 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_505 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_517 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_521 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_525 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_558 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_570 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_580 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_622 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_627 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_645 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_666 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_673 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_689 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_728 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_14 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_73 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_124 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_127 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_137 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_414 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_424 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_433 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_444 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_455 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_478 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_490 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_31_495 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_503 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_505 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_516 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_520 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_527 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_539 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_602 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_630 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_638 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_647 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_671 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_713 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_722 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_22 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_74 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_95 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_104 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_187 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_262 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_303 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_318 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_358 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_378 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_387 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_434 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_32_443 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_462 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_474 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_32_477 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_483 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_32_489 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_495 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_32_503 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_509 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_589 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_594 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_636 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_643 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_657 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_677 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_699 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_18 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_159 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_221 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_244 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_260 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_268 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_361 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_437 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_446 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_33_469 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_475 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_491 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_512 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_601 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_651 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_671 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_675 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_702 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_727 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_45 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_130 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_276 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_309 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_318 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_344 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_34_453 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_34_470 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_477 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_560 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_575 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_585 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_624 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_643 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_650 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_692 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_7 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_50 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_66 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_196 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_202 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_250 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_288 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_294 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_337 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_451 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_455 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_461 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_473 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_480 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_35_485 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_35_493 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_502 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_514 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_581 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_613 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_623 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_631 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_647 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_671 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_703 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_93 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_220 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_314 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_354 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_390 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_398 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_36_469 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_475 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_487 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_36_501 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_509 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_535 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_568 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_668 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_689 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_732 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_46 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_59 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_147 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_151 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_157 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_37_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_257 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_261 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_37_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_337 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_361 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_408 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_439 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_37_500 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_505 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_533 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_557 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_671 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_692 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_96 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_137 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_147 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_158 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_192 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_201 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_38_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_38_268 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_38_276 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_425 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_431 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_38_464 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_475 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_38_489 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_38_506 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_587 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_618 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_635 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_656 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_667 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_732 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_140 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_203 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_231 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_39_265 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_39_294 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_352 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_433 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_460 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_468 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_486 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_489 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_39_496 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_531 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_671 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_687 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_39 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_69 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_40_205 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_211 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_220 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_239 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_40_265 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_274 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_40_287 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_40_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_338 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_391 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_40_451 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_475 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_522 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_531 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_533 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_539 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_572 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_582 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_635 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_659 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_33 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_63 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_150 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_157 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_41_162 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_177 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_41_206 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_41_220 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_41_230 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_242 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_41_252 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_258 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_41_299 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_342 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_361 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_391 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_449 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_472 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_498 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_503 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_599 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_671 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_681 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_7 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_78 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_117 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_42_129 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_42_137 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_42_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_42_173 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_42_178 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_42_191 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_42_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_205 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_247 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_42_274 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_280 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_42_300 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_309 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_42_322 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_330 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_363 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_365 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_409 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_456 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_519 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_587 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_638 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_677 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_694 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_724 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_71 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_135 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_43_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_43_210 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_43_221 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_230 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_261 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_43_283 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_43_314 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_320 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_340 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_376 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_385 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_426 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_523 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_565 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_705 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_116 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_124 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_128 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_216 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_227 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_247 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_261 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_44_285 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_44_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_309 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_326 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_44_383 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_475 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_540 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_583 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_645 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_688 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_712 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_43 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_173 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_187 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_202 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_208 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_215 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_45_287 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_299 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_311 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_362 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_379 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_443 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_457 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_491 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_503 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_508 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_523 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_529 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_548 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_568 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_576 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_603 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_671 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_719 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_112 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_127 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_202 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_211 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_259 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_46_275 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_46_295 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_301 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_309 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_46_322 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_46_330 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_338 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_349 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_46_377 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_529 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_631 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_699 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_719 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_47 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_68 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_47_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_155 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_162 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_204 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_218 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_47_318 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_326 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_47_332 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_373 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_401 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_431 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_466 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_505 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_533 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_549 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_563 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_48_123 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_129 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_132 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_48_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_48_153 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_48_157 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_48_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_176 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_187 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_48_194 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_48_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_203 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_212 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_267 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_48_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_48_309 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_48_345 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_357 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_374 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_399 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_419 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_448 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_460 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_475 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_479 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_538 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_643 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_50 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_49_91 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_98 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_49_102 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_49_151 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_155 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_49_171 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_49_186 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_190 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_221 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_260 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_272 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_299 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_49_307 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_49_344 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_49_376 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_412 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_421 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_503 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_561 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_578 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_592 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_671 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_14 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_58 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_50_98 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_50_128 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_50_150 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_154 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_50_157 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_50_180 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_201 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_215 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_236 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_290 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_50_301 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_50_314 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_50_321 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_327 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_342 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_50_347 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_359 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_373 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_421 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_466 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_475 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_496 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_502 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_526 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_597 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_611 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_633 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_699 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_51_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_61 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_51_65 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_69 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_51_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_51_106 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_51_132 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_155 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_181 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_198 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_230 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_260 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_269 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_51_304 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_51_313 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_317 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_51_320 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_326 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_337 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_51_356 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_379 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_385 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_449 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_480 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_539 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_577 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_696 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_36 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_61 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_52_71 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_52_97 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_123 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_52_135 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_168 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_52_178 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_203 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_259 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_306 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_309 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_327 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_337 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_346 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_52_365 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_52_386 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_400 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_411 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_445 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_454 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_533 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_567 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_678 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_53_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_87 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_53_96 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_53_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_153 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_200 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_53_211 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_230 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_258 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_275 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_298 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_53_307 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_53_317 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_323 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_329 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_337 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_53_342 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_350 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_53_385 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_391 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_393 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_418 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_428 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_434 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_512 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_559 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_628 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_19 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_93 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_109 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_126 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_54_129 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_54_137 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_153 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_54_165 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_54_179 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_183 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_54_190 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_54_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_54_205 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_54_303 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_330 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_337 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_353 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_363 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_54_367 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_373 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_379 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_387 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_423 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_432 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_440 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_475 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_531 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_533 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_587 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_643 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_686 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_59 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_55_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_84 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_96 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_55_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_119 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_130 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_55_156 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_55_178 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_192 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_204 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_212 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_218 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_233 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_286 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_308 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_351 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_372 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_376 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_55_401 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_405 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_412 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_498 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_615 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_617 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_627 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_693 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_707 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_56_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_56_119 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_56_131 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_56_148 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_160 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_56_164 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_172 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_199 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_56_205 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_322 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_328 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_365 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_387 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_411 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_469 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_587 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_643 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_674 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_57_87 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_57_99 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_57_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_57_128 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_134 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_57_150 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_176 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_204 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_214 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_262 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_308 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_322 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_356 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_447 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_467 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_578 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_610 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_56 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_58_63 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_75 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_58_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_91 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_100 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_58_109 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_115 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_58_125 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_58_137 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_58_144 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_205 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_58_215 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_58_227 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_235 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_309 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_371 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_475 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_531 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_655 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_694 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_709 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_732 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_19 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_47 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_59_78 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_86 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_59_107 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_59_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_59_130 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_59_171 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_198 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_59_216 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_232 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_238 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_259 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_286 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_328 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_484 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_559 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_570 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_34 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_60_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_60_92 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_60_99 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_60_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_137 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_154 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_60_172 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_60_180 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_199 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_60_213 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_240 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_249 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_432 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_475 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_493 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_662 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_732 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_61_101 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_109 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_61_132 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_203 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_221 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_228 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_454 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_519 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_559 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_587 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_615 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_671 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_61_673 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_701 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_11 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_19 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_40 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_61 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_62_70 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_62_78 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_62_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_116 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_126 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_178 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_202 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_62_234 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_255 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_331 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_365 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_379 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_419 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_450 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_475 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_495 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_533 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_612 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_633 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_643 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_692 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_48 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_63_62 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_63_68 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_97 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_63_116 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_134 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_154 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_63_199 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_63_235 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_245 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_252 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_291 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_337 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_366 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_419 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_428 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_496 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_662 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_64_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_101 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_64_125 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_154 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_64_180 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_184 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_64_201 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_64_209 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_64_219 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_64_231 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_64_239 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_298 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_419 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_469 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_501 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_514 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_526 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_533 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_587 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_619 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_64_634 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_723 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_732 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_65_46 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_65_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_65_74 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_65_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_65_91 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_174 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_65_182 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_65_201 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_65_219 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_65_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_294 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_342 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_399 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_487 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_597 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_639 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_699 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_66_36 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_66_45 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_66_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_66_92 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_66_100 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_66_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_120 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_66_194 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_66_203 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_66_211 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_66_230 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_234 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_66_237 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_294 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_307 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_373 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_393 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_406 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_467 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_475 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_519 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_531 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_591 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_618 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_659 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_688 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_699 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_710 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_720 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_67_35 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_67_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_67_109 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_67_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_150 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_67_153 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_67_166 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_67_176 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_180 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_67_239 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_67_248 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_67_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_67_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_285 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_323 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_67_333 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_337 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_563 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_671 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_686 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_5 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_68_10 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_18 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_32 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_38 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_60 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_64 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_68_68 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_68_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_97 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_68_107 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_115 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_68_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_68_168 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_68_180 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_68_192 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_68_201 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_68_213 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_68_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_68_231 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_237 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_68_246 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_307 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_363 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_68_365 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_369 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_389 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_465 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_477 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_498 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_597 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_638 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_699 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_69_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_69_43 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_64 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_75 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_69_107 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_69_135 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_69_148 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_69_185 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_69_206 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_214 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_69_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_69_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_294 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_347 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_391 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_407 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_447 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_494 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_503 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_573 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_622 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_671 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_686 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_719 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_37 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_60 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_70_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_70_100 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_104 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_70_128 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_173 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_179 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_70_191 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_70_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_217 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_229 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_70_241 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_260 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_266 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_292 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_70_295 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_311 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_70_321 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_70_356 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_368 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_399 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_414 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_475 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_577 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_606 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_699 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_71_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_71_16 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_22 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_65 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_71_71 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_71_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_71_88 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_71_118 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_126 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_135 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_140 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_71_149 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_166 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_192 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_197 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_209 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_71_219 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_228 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_71_238 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_266 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_286 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_329 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_71_333 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_71_361 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_365 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_71_372 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_376 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_71_384 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_422 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_503 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_536 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_546 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_561 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_617 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_666 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_10 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_72_18 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_72_36 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_42 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_72_70 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_72_81 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_72_146 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_152 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_72_160 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_72_180 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_209 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_72_221 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_302 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_72_337 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_382 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_477 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_505 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_546 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_638 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_660 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_26 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_73_38 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_42 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_73_86 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_118 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_73_155 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_180 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_207 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_73_219 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_73_235 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_284 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_315 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_335 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_73_385 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_389 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_435 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_487 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_509 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_559 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_600 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_617 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_699 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_74_19 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_58 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_74_79 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_127 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_74_130 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_141 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_74_153 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_74_184 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_74_242 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_298 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_309 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_336 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_74_361 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_365 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_448 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_457 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_475 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_494 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_540 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_550 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_570 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_580 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_594 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_643 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_683 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_10 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_17 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_25 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_75_46 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_50 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_75_65 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_73 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_120 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_132 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_75_144 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_180 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_183 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_75_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_235 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_75_244 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_252 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_292 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_304 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_316 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_75_323 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_327 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_75_333 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_75_339 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_345 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_351 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_75_354 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_75_382 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_422 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_458 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_462 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_535 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_589 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_617 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_693 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_76_45 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_76_56 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_76_73 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_76_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_120 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_148 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_181 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_76_239 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_245 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_317 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_411 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_463 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_475 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_547 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_647 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_708 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_732 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_46 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_84 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_77_150 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_176 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_219 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_238 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_275 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_407 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_484 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_608 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_626 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_698 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_78_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_10 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_78_34 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_72 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_78_130 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_78_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_78_159 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_78_175 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_78_219 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_78_229 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_255 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_78_278 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_282 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_287 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_318 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_383 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_419 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_444 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_454 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_540 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_667 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_79_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_13 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_79_25 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_31 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_79_44 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_158 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_79_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_79_202 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_79_236 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_242 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_252 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_264 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_79_275 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_295 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_335 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_433 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_443 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_512 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_528 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_561 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_570 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_619 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_79_693 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_6 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_13 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_80_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_70 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_80_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_94 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_120 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_132 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_159 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_199 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_80_213 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_80_235 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_80_250 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_80_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_268 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_80_304 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_343 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_80_391 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_446 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_456 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_488 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_526 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_533 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_543 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_568 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_608 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_617 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_628 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_671 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_699 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_708 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_81_30 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_81_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_81_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_81_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_81_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_81_137 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_81_145 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_81_155 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_81_211 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_81_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_81_277 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_81_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_81_291 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_81_299 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_81_354 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_81_451 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_81_472 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_81_505 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_81_534 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_81_576 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_81_658 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_81_675 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_82_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_82_62 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_82_153 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_82_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_82_177 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_82_186 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_82_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_82_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_82_205 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_82_209 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_82_215 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_82_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_82_233 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_82_257 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_82_282 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_82_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_82_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_82_303 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_82_320 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_82_347 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_82_361 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_82_419 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_82_435 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_82_470 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_82_560 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_82_681 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_82_699 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_82_715 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_82_732 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_83_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_83_37 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_83_46 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_83_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_83_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_83_137 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_83_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_83_151 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_83_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_83_210 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_83_222 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_83_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_83_239 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_83_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_83_288 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_83_295 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_83_337 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_83_349 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_83_381 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_83_449 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_83_527 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_83_573 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_83_617 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_83_666 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_83_681 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_84_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_84_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_84_87 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_84_112 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_84_119 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_84_127 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_84_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_84_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_84_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_84_265 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_84_374 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_84_606 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_84_643 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_84_692 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_85_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_85_48 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_85_59 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_85_70 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_85_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_85_129 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_85_158 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_85_166 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_85_186 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_85_206 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_85_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_85_267 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_85_337 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_85_382 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_85_418 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_85_427 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_85_451 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_85_513 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_85_581 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_85_634 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_85_700 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_86_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_86_69 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_86_122 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_86_152 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_86_156 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_86_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_86_205 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_86_218 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_86_230 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_86_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_86_260 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_86_278 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_86_338 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_86_344 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_86_353 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_86_399 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_86_459 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_86_488 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_86_579 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_86_632 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_86_643 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_86_651 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_86_678 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_87_14 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_87_35 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_87_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_87_70 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_87_81 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_87_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_87_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_87_137 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_87_148 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_87_156 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_87_174 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_87_200 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_87_222 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_87_245 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_87_252 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_87_260 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_87_286 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_87_307 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_87_391 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_87_439 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_87_553 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_87_571 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_87_619 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_87_678 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_87_719 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_88_32 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_88_50 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_88_128 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_88_134 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_88_143 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_88_154 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_88_162 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_88_166 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_88_170 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_88_217 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_88_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_88_229 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_88_267 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_88_340 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_88_429 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_88_511 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_88_547 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_88_616 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_88_647 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_88_684 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_88_712 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_89_69 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_89_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_89_97 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_89_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_89_175 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_89_187 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_89_198 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_89_202 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_89_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_89_233 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_89_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_89_290 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_89_378 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_89_397 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_89_538 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_89_590 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_89_628 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_89_671 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_89_683 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_90_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_90_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_90_36 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_90_66 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_90_78 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_90_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_90_118 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_90_132 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_90_190 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_90_205 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_90_211 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_90_220 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_90_224 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_90_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_90_367 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_90_477 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_90_510 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_90_566 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_90_598 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_90_622 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_90_645 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_90_690 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_90_699 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_90_732 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_91_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_91_84 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_91_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_91_178 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_91_187 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_91_209 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_91_229 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_91_328 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_91_352 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_91_413 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_91_420 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_91_547 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_91_568 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_91_594 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_91_653 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_91_675 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_91_698 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_92_20 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_92_46 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_92_175 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_92_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_92_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_92_201 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_92_221 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_92_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_92_246 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_92_392 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_92_414 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_92_427 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_92_479 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_92_537 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_92_547 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_92_617 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_92_628 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_92_715 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_93_48 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_93_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_93_68 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_93_120 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_93_129 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_93_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_93_149 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_93_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_93_176 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_93_188 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_93_199 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_93_217 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_93_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_93_342 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_93_395 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_93_436 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_93_462 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_93_485 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_93_561 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_93_605 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_93_690 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_93_701 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_94_120 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_94_129 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_94_155 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_94_164 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_94_178 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_94_191 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_94_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_94_231 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_94_242 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_94_335 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_94_342 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_94_359 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_94_382 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_94_458 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_94_525 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_94_547 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_94_569 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_94_583 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_94_591 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_94_623 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_94_675 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_94_697 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_94_712 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_95_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_95_62 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_95_115 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_95_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_95_154 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_95_162 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_95_197 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_95_209 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_95_229 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_95_315 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_95_337 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_95_367 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_95_380 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_95_432 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_95_525 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_95_624 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_95_671 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_96_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_96_43 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_96_90 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_96_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_96_149 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_96_172 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_96_186 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_96_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_96_201 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_96_216 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_96_220 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_96_230 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_96_239 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_96_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_96_270 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_96_287 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_96_314 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_96_317 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_96_365 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_96_401 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_96_407 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_96_414 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_96_471 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_96_482 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_96_574 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_96_690 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_96_712 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_97_41 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_97_53 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_97_68 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_97_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_97_127 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_97_158 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_97_166 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_97_175 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_97_187 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_97_200 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_97_208 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_97_219 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_97_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_97_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_97_357 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_97_542 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_97_619 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_97_651 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_98_33 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_98_39 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_98_47 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_98_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_98_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_98_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_98_158 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_98_260 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_98_294 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_98_352 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_98_428 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_98_495 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_98_637 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_98_666 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_98_699 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_98_701 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_98_732 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_99_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_99_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_99_118 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_99_125 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_99_129 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_99_155 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_99_159 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_99_162 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_99_173 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_99_183 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_99_201 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_99_228 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_99_244 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_99_308 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_99_515 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_99_556 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_99_631 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_99_732 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_100_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_100_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_100_62 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_100_78 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_100_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_100_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_100_134 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_100_146 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_100_160 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_100_171 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_100_367 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_100_401 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_100_423 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_100_549 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_100_643 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_100_724 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_101_11 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_101_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_101_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_101_81 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_101_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_101_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_101_119 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_101_125 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_101_129 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_101_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_101_324 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_101_399 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_101_427 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_101_464 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_101_494 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_101_557 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_101_651 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_102_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_102_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_102_46 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_102_120 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_102_132 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_102_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_102_210 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_102_230 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_102_246 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_102_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_102_301 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_102_355 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_102_382 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_102_404 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_102_419 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_102_459 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_102_574 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_102_712 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_103_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_103_10 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_103_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_103_64 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_103_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_103_106 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_103_120 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_103_162 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_103_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_103_221 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_103_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_103_257 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_103_287 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_103_327 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_103_374 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_103_445 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_103_530 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_103_579 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_104_14 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_104_19 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_104_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_104_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_104_38 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_104_50 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_104_62 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_104_72 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_104_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_104_99 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_104_116 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_104_150 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_104_183 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_104_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_104_215 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_104_219 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_104_245 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_104_267 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_104_303 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_104_363 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_104_408 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_104_465 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_104_495 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_104_547 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_104_559 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_104_666 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_104_689 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_105_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_105_62 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_105_94 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_105_102 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_105_126 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_105_131 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_105_140 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_105_187 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_105_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_105_205 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_105_210 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_105_214 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_105_222 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_105_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_105_333 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_105_352 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_105_391 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_105_399 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_105_443 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_105_462 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_105_491 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_105_519 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_105_559 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_105_578 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_105_659 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_105_681 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_105_711 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_106_37 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_106_66 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_106_93 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_106_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_106_144 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_106_153 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_106_177 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_106_182 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_106_194 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_106_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_106_247 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_106_300 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_106_307 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_106_320 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_106_358 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_106_399 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_106_451 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_106_477 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_106_520 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_106_610 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_106_626 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_106_645 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_107_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_107_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_107_90 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_107_99 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_107_116 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_107_145 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_107_160 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_107_183 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_107_191 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_107_222 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_107_230 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_107_315 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_107_322 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_107_368 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_107_377 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_107_389 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_107_393 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_107_428 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_107_449 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_107_501 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_107_591 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_107_615 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_107_642 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_107_651 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_108_44 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_108_52 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_108_64 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_108_71 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_108_81 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_108_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_108_95 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_108_99 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_108_123 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_108_146 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_108_167 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_108_179 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_108_194 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_108_230 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_108_244 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_108_266 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_108_294 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_108_342 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_108_367 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_108_388 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_108_394 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_108_402 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_108_406 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_108_411 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_108_419 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_108_421 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_108_457 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_108_486 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_108_556 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_108_563 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_108_589 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_108_674 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_108_699 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_109_23 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_109_35 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_109_70 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_109_92 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_109_100 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_109_118 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_109_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_109_154 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_109_165 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_109_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_109_173 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_109_199 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_109_213 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_109_222 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_109_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_109_232 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_109_236 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_109_263 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_109_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_109_337 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_109_382 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_109_404 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_109_430 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_109_486 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_110_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_110_102 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_110_107 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_110_119 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_110_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_110_144 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_110_177 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_110_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_110_226 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_110_235 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_110_249 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_110_401 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_110_405 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_110_416 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_110_425 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_110_431 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_110_473 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_110_531 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_110_587 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_110_596 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_110_617 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_110_628 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_110_661 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_110_722 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_111_50 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_111_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_111_68 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_111_92 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_111_98 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_111_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_111_118 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_111_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_111_165 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_111_205 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_111_277 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_111_356 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_111_362 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_111_365 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_111_369 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_111_381 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_111_389 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_111_402 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_111_424 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_111_451 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_111_460 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_111_536 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_111_559 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_111_570 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_111_619 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_111_675 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_111_700 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_112_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_112_32 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_112_65 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_112_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_112_81 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_112_92 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_112_157 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_112_174 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_112_232 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_112_241 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_112_292 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_112_363 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_112_375 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_112_383 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_112_403 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_112_440 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_112_452 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_112_494 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_112_529 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_112_550 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_112_587 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_112_598 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_112_643 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_112_647 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_112_699 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_112_732 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_113_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_113_65 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_113_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_113_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_113_122 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_113_132 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_113_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_113_140 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_113_147 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_113_156 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_113_164 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_113_192 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_113_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_113_233 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_113_241 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_113_266 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_113_278 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_113_292 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_113_335 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_113_337 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_113_348 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_113_369 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_113_390 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_113_449 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_113_485 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_113_497 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_113_505 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_113_559 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_113_566 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_113_625 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_113_662 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_113_691 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_114_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_114_19 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_114_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_114_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_114_37 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_114_43 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_114_70 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_114_81 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_114_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_114_146 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_114_175 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_114_186 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_114_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_114_212 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_114_230 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_114_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_114_261 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_114_273 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_114_287 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_114_295 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_114_363 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_114_365 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_114_369 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_114_378 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_114_382 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_114_430 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_114_477 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_114_546 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_114_611 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_114_643 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_114_688 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_114_699 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_114_732 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_115_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_115_10 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_115_22 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_115_34 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_115_60 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_115_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_115_93 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_115_102 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_115_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_115_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_115_135 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_115_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_115_192 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_115_215 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_115_234 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_115_246 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_115_260 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_115_272 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_115_291 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_115_319 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_115_352 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_115_379 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_115_446 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_115_546 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_115_551 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_115_582 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_115_661 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_115_719 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_116_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_116_17 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_116_25 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_116_29 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_116_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_116_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_116_94 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_116_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_116_149 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_116_160 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_116_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_116_176 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_116_194 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_116_202 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_116_216 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_116_243 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_116_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_116_253 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_116_265 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_116_275 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_116_287 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_116_299 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_116_303 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_116_326 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_116_363 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_116_376 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_116_438 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_116_446 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_116_564 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_116_585 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_116_596 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_116_653 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_116_688 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_116_699 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_116_722 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_117_28 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_117_40 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_117_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_117_59 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_117_63 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_117_69 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_117_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_117_166 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_117_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_117_188 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_117_236 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_117_260 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_117_268 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_117_274 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_117_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_117_295 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_117_354 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_117_388 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_117_393 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_117_408 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_117_543 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_117_595 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_117_661 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_118_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_118_12 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_118_33 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_118_39 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_118_46 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_118_53 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_118_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_118_97 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_118_119 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_118_151 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_118_172 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_118_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_118_260 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_118_282 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_118_286 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_118_309 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_118_320 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_118_419 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_118_442 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_118_473 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_118_533 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_118_547 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_118_597 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_118_604 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_118_613 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_118_621 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_118_626 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_118_643 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_118_672 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_118_705 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_118_711 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_118_732 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_119_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_119_35 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_119_42 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_119_49 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_119_53 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_119_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_119_65 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_119_73 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_119_79 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_119_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_119_85 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_119_97 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_119_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_119_188 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_119_205 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_119_212 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_119_218 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_119_221 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_119_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_119_229 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_119_235 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_119_247 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_119_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_119_253 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_119_265 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_119_277 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_119_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_119_287 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_119_307 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_119_393 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_119_397 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_119_403 (.VPWR(vccd1),
    .VGND(vssd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_119_415 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_119_419 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_119_429 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_119_437 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_119_449 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_119_464 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_119_501 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_119_533 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_119_569 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_119_584 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_119_587 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_119_593 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_119_602 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_119_613 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_119_617 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_119_636 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_119_643 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_119_649 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_119_660 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_119_673 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_119_684 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
endmodule
