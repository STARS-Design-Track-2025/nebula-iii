`default_nettype none
/////////////////////////////////////////////////////////////////
// HEADER 
//
// Module : t01_clkdiv1hz
// Description : takes 25mhz clock and turns it into 1 hz enable
// 
//
/////////////////////////////////////////////////////////////////
module t01_clkdiv1hz (
    input logic clk, rst, //25mhz -> 1hz
    input logic [24:0] scoremod,
    input logic speed_up,
    input logic [1:0] top_level_state, 
    output logic newclk
);

    logic [25:0] count, count_n;
    logic newclk_n;
    logic [25:0] threshold, clk_speed_div; 

    // assign the clk speed based on Tetris game mode 
    assign clk_speed_div = top_level_state == 2'b01 ? 26'd1_250_000 : 26'd100; 

    always_ff @(posedge clk, posedge rst) begin
       if (rst) begin
            count <= '0;
            newclk <= '0;
       end else begin
            count <= count_n;
            newclk <= newclk_n;
       end
    end

    always_comb begin
        count_n = count;
        newclk_n = '1;
        threshold = speed_up ? clk_speed_div : 26'd12_500_000 - scoremod; // clock adjustment 
        if (count < threshold) begin // updated to half a huzz
            count_n = count + 1;
        end else begin
            count_n = '0;
            newclk_n = '0;
        end
    end
endmodule