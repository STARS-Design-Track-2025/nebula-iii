* NGSPICE file created from team_00.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_4 abstract view
.subckt sky130_fd_sc_hd__fill_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_40_12 abstract view
.subckt sky130_ef_sc_hd__decap_40_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_8 abstract view
.subckt sky130_fd_sc_hd__fill_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufinv_16 abstract view
.subckt sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

.subckt team_00 clk done en gpio_in[0] gpio_in[10] gpio_in[11] gpio_in[12] gpio_in[13]
+ gpio_in[14] gpio_in[15] gpio_in[16] gpio_in[17] gpio_in[18] gpio_in[19] gpio_in[1]
+ gpio_in[20] gpio_in[21] gpio_in[22] gpio_in[23] gpio_in[24] gpio_in[25] gpio_in[26]
+ gpio_in[27] gpio_in[28] gpio_in[29] gpio_in[2] gpio_in[30] gpio_in[31] gpio_in[32]
+ gpio_in[33] gpio_in[3] gpio_in[4] gpio_in[5] gpio_in[6] gpio_in[7] gpio_in[8] gpio_in[9]
+ gpio_oeb[0] gpio_oeb[10] gpio_oeb[11] gpio_oeb[12] gpio_oeb[13] gpio_oeb[14] gpio_oeb[15]
+ gpio_oeb[16] gpio_oeb[17] gpio_oeb[18] gpio_oeb[19] gpio_oeb[1] gpio_oeb[20] gpio_oeb[21]
+ gpio_oeb[22] gpio_oeb[23] gpio_oeb[24] gpio_oeb[25] gpio_oeb[26] gpio_oeb[27] gpio_oeb[28]
+ gpio_oeb[29] gpio_oeb[2] gpio_oeb[30] gpio_oeb[31] gpio_oeb[32] gpio_oeb[33] gpio_oeb[3]
+ gpio_oeb[4] gpio_oeb[5] gpio_oeb[6] gpio_oeb[7] gpio_oeb[8] gpio_oeb[9] gpio_out[0]
+ gpio_out[10] gpio_out[11] gpio_out[12] gpio_out[13] gpio_out[14] gpio_out[15] gpio_out[16]
+ gpio_out[17] gpio_out[18] gpio_out[19] gpio_out[1] gpio_out[20] gpio_out[21] gpio_out[22]
+ gpio_out[23] gpio_out[24] gpio_out[25] gpio_out[26] gpio_out[27] gpio_out[28] gpio_out[29]
+ gpio_out[2] gpio_out[30] gpio_out[31] gpio_out[32] gpio_out[33] gpio_out[3] gpio_out[4]
+ gpio_out[5] gpio_out[6] gpio_out[7] gpio_out[8] gpio_out[9] la_data_in[0] la_data_in[10]
+ la_data_in[11] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16]
+ la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20] la_data_in[21]
+ la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26] la_data_in[27]
+ la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31] la_data_in[3]
+ la_data_in[4] la_data_in[5] la_data_in[6] la_data_in[7] la_data_in[8] la_data_in[9]
+ la_data_out[0] la_data_out[10] la_data_out[11] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24]
+ la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29]
+ la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[3] la_data_out[4] la_data_out[5]
+ la_data_out[6] la_data_out[7] la_data_out[8] la_data_out[9] la_oenb[0] la_oenb[10]
+ la_oenb[11] la_oenb[12] la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17]
+ la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23]
+ la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2]
+ la_oenb[30] la_oenb[31] la_oenb[3] la_oenb[4] la_oenb[5] la_oenb[6] la_oenb[7] la_oenb[8]
+ la_oenb[9] nrst prescaler[0] prescaler[10] prescaler[11] prescaler[12] prescaler[13]
+ prescaler[1] prescaler[2] prescaler[3] prescaler[4] prescaler[5] prescaler[6] prescaler[7]
+ prescaler[8] prescaler[9] vccd1 vssd1
XFILLER_79_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_94_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_27_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_39_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_67_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_82_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_35_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_22_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_52_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_50_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__0703__A net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_58_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_85_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_73_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_93_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_26_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_14_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_9_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_41_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__0613__A net18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1270_ _0581_ _0591_ _0604_ vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__and3_1
XFILLER_95_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_76_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_49_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_47_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_64_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_19_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_17_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_32_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0985_ net13 _0019_ _0373_ _0374_ vssd1 vssd1 vccd1 vccd1 _0375_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_74_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_87_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout116 net117 vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__clkbuf_2
Xfanout105 count\[2\] vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__clkbuf_2
XFILLER_101_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_67_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_55_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xteam_00_148 vssd1 vssd1 vccd1 vccd1 team_00_148/HI la_data_out[22] sky130_fd_sc_hd__conb_1
Xteam_00_137 vssd1 vssd1 vccd1 vccd1 team_00_137/HI la_data_out[11] sky130_fd_sc_hd__conb_1
Xteam_00_126 vssd1 vssd1 vccd1 vccd1 team_00_126/HI la_data_out[0] sky130_fd_sc_hd__conb_1
XFILLER_27_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_63_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_12_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_2_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_77_147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_46_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_92_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_33_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__0608__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_61_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_53_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_52_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0770_ _0152_ _0159_ _0158_ vssd1 vssd1 vccd1 vccd1 _0160_ sky130_fd_sc_hd__a21o_1
XFILLER_96_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_69_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_96_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1253_ _0577_ _0599_ vssd1 vssd1 vccd1 vccd1 _0600_ sky130_fd_sc_hd__and2_1
XFILLER_56_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1317__RESET_B net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1184_ _0186_ clk_divider.next_count\[13\] vssd1 vssd1 vccd1 vccd1 _0542_ sky130_fd_sc_hd__xnor2_1
XFILLER_91_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_20_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_60_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_20_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0968_ clk_divider.count_out\[15\] _0182_ vssd1 vssd1 vccd1 vccd1 _0358_ sky130_fd_sc_hd__nand2_1
XFILLER_20_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0899_ _0281_ _0278_ vssd1 vssd1 vccd1 vccd1 _0289_ sky130_fd_sc_hd__nand2b_1
XFILLER_99_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__0700__B net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_59_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_28_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_15_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_28_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_83_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_43_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_30_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_70_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_23_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_11_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_7_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_21_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_94_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_78_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_2_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_78_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_38_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_78_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1281__X net81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_29_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_61_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0822_ _0203_ _0205_ _0206_ vssd1 vssd1 vccd1 vccd1 _0212_ sky130_fd_sc_hd__o21bai_1
X_0753_ _0140_ _0141_ vssd1 vssd1 vccd1 vccd1 _0143_ sky130_fd_sc_hd__xnor2_1
X_0684_ net16 net15 vssd1 vssd1 vccd1 vccd1 _0074_ sky130_fd_sc_hd__xor2_1
XFILLER_50_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_88_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_71_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1305_ clknet_2_1__leaf_clk clk_divider.next_count\[21\] net121 vssd1 vssd1 vccd1
+ vccd1 clk_divider.count_out\[21\] sky130_fd_sc_hd__dfrtp_1
X_1236_ _0000_ _0588_ _0590_ vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__and3_1
X_1167_ clk_divider.count_out\[25\] net109 _0524_ _0527_ net98 vssd1 vssd1 vccd1 vccd1
+ clk_divider.next_count\[25\] sky130_fd_sc_hd__o221a_1
XFILLER_52_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_25_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_52_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1098_ clk_divider.count_out\[14\] _0465_ vssd1 vssd1 vccd1 vccd1 _0470_ sky130_fd_sc_hd__xor2_1
XFILLER_40_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_20_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_60_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1315__CLK clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_55_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_26_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_24_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_31_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_34_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_43_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1021__A2 _0199_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_3_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_78_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_78_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_93_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_75_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1021_ net113 _0199_ _0027_ vssd1 vssd1 vccd1 vccd1 _0410_ sky130_fd_sc_hd__a21oi_1
XFILLER_34_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_34_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_98_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_22_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_61_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_32_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0805_ _0169_ _0194_ vssd1 vssd1 vccd1 vccd1 _0195_ sky130_fd_sc_hd__or2_2
X_0736_ net13 _0105_ vssd1 vssd1 vccd1 vccd1 _0126_ sky130_fd_sc_hd__xnor2_1
XFILLER_89_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0667_ _0047_ _0055_ vssd1 vssd1 vccd1 vccd1 _0057_ sky130_fd_sc_hd__xnor2_2
XFILLER_97_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_84_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_68_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_44_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1219_ _0549_ _0562_ _0576_ vssd1 vssd1 vccd1 vccd1 clk_divider.next_flag sky130_fd_sc_hd__nor3_1
XFILLER_37_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_80_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_91_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_0_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_75_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input18_A prescaler[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_16_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_16_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_45_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__0616__A net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_16_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_100_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_8_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_8_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_100_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_79_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1182__A _0199_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_94_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_65_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_37_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1004_ _0344_ _0393_ _0336_ _0340_ vssd1 vssd1 vccd1 vccd1 _0394_ sky130_fd_sc_hd__o211a_1
XFILLER_62_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_50_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_34_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_77_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0719_ _0010_ _0011_ vssd1 vssd1 vccd1 vccd1 _0109_ sky130_fd_sc_hd__nor2_1
XFILLER_17_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_88_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_13_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_40_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0983__A1 net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput31 net31 vssd1 vssd1 vccd1 vccd1 gpio_oeb[18] sky130_fd_sc_hd__buf_2
Xoutput42 net42 vssd1 vssd1 vccd1 vccd1 gpio_oeb[28] sky130_fd_sc_hd__buf_2
Xoutput64 net64 vssd1 vssd1 vccd1 vccd1 gpio_out[17] sky130_fd_sc_hd__buf_2
Xoutput75 net75 vssd1 vssd1 vccd1 vccd1 gpio_out[27] sky130_fd_sc_hd__buf_2
Xoutput53 net53 vssd1 vssd1 vccd1 vccd1 gpio_oeb[7] sky130_fd_sc_hd__buf_2
XFILLER_95_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xoutput86 net86 vssd1 vssd1 vccd1 vccd1 gpio_out[6] sky130_fd_sc_hd__buf_2
XFILLER_48_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_62_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_32_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_86_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_27_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_82_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_35_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_50_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_89_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_77_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_93_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_85_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_58_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_26_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_26_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_53_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_9_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_42_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_11_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_97_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_95_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_3_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1163__C net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_64_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_19_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_83_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_32_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_80_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0984_ _0010_ clk_divider.count_out\[7\] vssd1 vssd1 vccd1 vccd1 _0374_ sky130_fd_sc_hd__nor2_1
XFILLER_8_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_74_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout106 count\[1\] vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__clkbuf_2
Xfanout117 net118 vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__clkbuf_2
XFILLER_86_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
Xteam_00_138 vssd1 vssd1 vccd1 vccd1 team_00_138/HI la_data_out[12] sky130_fd_sc_hd__conb_1
Xteam_00_149 vssd1 vssd1 vccd1 vccd1 team_00_149/HI la_data_out[23] sky130_fd_sc_hd__conb_1
Xteam_00_127 vssd1 vssd1 vccd1 vccd1 team_00_127/HI la_data_out[1] sky130_fd_sc_hd__conb_1
XFILLER_82_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_27_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_55_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_85_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_10_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1060__B1 _0036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_88_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_77_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_30 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_46_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_85_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_46_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_44_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_14_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_53_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_99_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_24_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_68_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1252_ net104 net106 net103 vssd1 vssd1 vccd1 vccd1 _0599_ sky130_fd_sc_hd__o21ai_1
XFILLER_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_64_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_37_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1183_ _0318_ _0518_ clk_divider.next_count\[2\] vssd1 vssd1 vccd1 vccd1 _0541_ sky130_fd_sc_hd__a21o_1
XFILLER_64_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_17_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_20_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0967_ clk_divider.count_out\[15\] _0182_ vssd1 vssd1 vccd1 vccd1 _0357_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_12_Right_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0898_ _0287_ vssd1 vssd1 vccd1 vccd1 _0288_ sky130_fd_sc_hd__inv_2
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_101_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_28_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_74_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_21_Right_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_82_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_23_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_7_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_21_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1033__B1 _0027_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_30_Right_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_94_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_fanout90_X net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_2_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_93_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_78_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_93_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_19_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_0_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_29_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_57_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0821_ _0049_ _0210_ _0209_ vssd1 vssd1 vccd1 vccd1 _0211_ sky130_fd_sc_hd__a21bo_1
X_0752_ _0140_ _0141_ vssd1 vssd1 vccd1 vccd1 _0142_ sky130_fd_sc_hd__nand2b_1
X_0683_ _0008_ _0009_ vssd1 vssd1 vccd1 vccd1 _0073_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_71_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_96_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1304_ clknet_2_1__leaf_clk clk_divider.next_count\[20\] net121 vssd1 vssd1 vccd1
+ vccd1 clk_divider.count_out\[20\] sky130_fd_sc_hd__dfrtp_1
XFILLER_96_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1235_ net105 _0023_ vssd1 vssd1 vccd1 vccd1 _0590_ sky130_fd_sc_hd__nor2_1
XFILLER_49_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_25_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1166_ net96 _0525_ _0526_ _0036_ vssd1 vssd1 vccd1 vccd1 _0527_ sky130_fd_sc_hd__a31o_1
XFILLER_52_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1097_ clk_divider.count_out\[14\] _0465_ vssd1 vssd1 vccd1 vccd1 _0469_ sky130_fd_sc_hd__and2_1
XFILLER_100_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_20_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_60_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1015__B1 _0199_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_75_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_75_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_28_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_90_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_28_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_26_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_34_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_11_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_7_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_50_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_59_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_6_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1020_ net97 _0408_ vssd1 vssd1 vccd1 vccd1 _0409_ sky130_fd_sc_hd__nand2_1
XFILLER_34_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_91_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_32_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0804_ _0167_ _0168_ vssd1 vssd1 vccd1 vccd1 _0194_ sky130_fd_sc_hd__and2_1
XFILLER_30_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0735_ _0122_ _0124_ vssd1 vssd1 vccd1 vccd1 _0125_ sky130_fd_sc_hd__nand2_1
X_0666_ _0047_ _0055_ vssd1 vssd1 vccd1 vccd1 _0056_ sky130_fd_sc_hd__nand2_1
XFILLER_69_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_69_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_97_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_57_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_57_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_72_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1218_ _0566_ _0570_ _0573_ _0575_ vssd1 vssd1 vccd1 vccd1 _0576_ sky130_fd_sc_hd__or4_1
XANTENNA__1301__RESET_B net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_9_Left_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1149_ _0508_ _0511_ _0512_ net98 vssd1 vssd1 vccd1 vccd1 clk_divider.next_count\[22\]
+ sky130_fd_sc_hd__o211a_1
XANTENNA__0706__B net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_21_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__0722__A net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_96_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_0_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout98_A net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_75_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1272__B _0605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_16_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_31_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_43_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_100_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_8_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_12_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_8_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_61_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_79_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_79_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_39_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_94_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_86_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_66_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1003_ _0348_ _0389_ _0390_ _0392_ vssd1 vssd1 vccd1 vccd1 _0393_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_37_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_22_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1305__CLK clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_6_Right_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_77_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0718_ _0106_ _0107_ vssd1 vssd1 vccd1 vccd1 _0108_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout100_A net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_89_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0649_ net8 _0038_ vssd1 vssd1 vccd1 vccd1 _0039_ sky130_fd_sc_hd__nand2_1
XFILLER_97_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_57_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0717__A net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_13_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_25_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_80_271 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_21_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1294__RESET_B net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput21 net21 vssd1 vssd1 vccd1 vccd1 done sky130_fd_sc_hd__buf_2
Xoutput43 net43 vssd1 vssd1 vccd1 vccd1 gpio_oeb[29] sky130_fd_sc_hd__buf_2
Xoutput32 net32 vssd1 vssd1 vccd1 vccd1 gpio_oeb[19] sky130_fd_sc_hd__buf_2
Xoutput65 net65 vssd1 vssd1 vccd1 vccd1 gpio_out[18] sky130_fd_sc_hd__buf_2
Xoutput76 net76 vssd1 vssd1 vccd1 vccd1 gpio_out[28] sky130_fd_sc_hd__buf_2
Xoutput54 net54 vssd1 vssd1 vccd1 vccd1 gpio_oeb[8] sky130_fd_sc_hd__buf_2
XFILLER_0_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
Xoutput87 net87 vssd1 vssd1 vccd1 vccd1 gpio_out[7] sky130_fd_sc_hd__buf_2
XFILLER_76_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_0_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_91_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_36_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_16_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_72_50 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_31_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_72_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_59_Right_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0726__A2 net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_79_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_68_Right_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_35_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_35_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_50_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_99_Left_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_77_Right_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1368__A net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_2_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_86_Right_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_93_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_85_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_73_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_45_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_26_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_95_Right_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_53_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_42_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_11_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__0708__A2 net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_1_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_3_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_95_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_76_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_91_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_19_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_47_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_83_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_32_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0983_ net13 _0019_ _0372_ vssd1 vssd1 vccd1 vccd1 _0373_ sky130_fd_sc_hd__o21ai_1
XFILLER_32_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_74_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout107 count\[0\] vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__clkbuf_2
Xfanout118 net48 vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__clkbuf_2
XFILLER_101_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_79_190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
Xteam_00_139 vssd1 vssd1 vccd1 vccd1 team_00_139/HI la_data_out[13] sky130_fd_sc_hd__conb_1
Xteam_00_128 vssd1 vssd1 vccd1 vccd1 team_00_128/HI la_data_out[2] sky130_fd_sc_hd__conb_1
XFILLER_67_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_27_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_55_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_27_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_85_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_11_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_6_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_37_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_46_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_58_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_18_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_61_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_14_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_99_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_53_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1174__C net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_96_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1251_ _0589_ _0598_ vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__nor2_1
XFILLER_76_160 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_37_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1182_ _0199_ clk_divider.next_count\[0\] clk_divider.next_count\[1\] vssd1 vssd1
+ vccd1 vccd1 _0540_ sky130_fd_sc_hd__or3_1
XFILLER_94_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_49_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_64_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_17_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_20_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_0966_ _0353_ _0354_ vssd1 vssd1 vccd1 vccd1 _0356_ sky130_fd_sc_hd__nand2_1
X_0897_ _0231_ _0264_ vssd1 vssd1 vccd1 vccd1 _0287_ sky130_fd_sc_hd__or2_1
XFILLER_87_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_67_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_27_Left_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_55_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_43_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_51_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_21_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_36_Left_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_94_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_78_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_48_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_93_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_19_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_45_Left_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_46_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_48_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_29_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_51 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_46_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__0635__A net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0820_ _0202_ _0208_ vssd1 vssd1 vccd1 vccd1 _0210_ sky130_fd_sc_hd__xor2_2
XPHY_EDGE_ROW_54_Left_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0751_ _0109_ _0119_ vssd1 vssd1 vccd1 vccd1 _0141_ sky130_fd_sc_hd__xnor2_1
X_0682_ _0045_ _0046_ vssd1 vssd1 vccd1 vccd1 _0072_ sky130_fd_sc_hd__xnor2_1
XFILLER_6_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_71_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_96_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_69_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1303_ clknet_2_1__leaf_clk clk_divider.next_count\[19\] net120 vssd1 vssd1 vccd1
+ vccd1 clk_divider.count_out\[19\] sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_63_Left_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_96_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_84_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1234_ _0585_ _0587_ vssd1 vssd1 vccd1 vccd1 _0589_ sky130_fd_sc_hd__or2_2
XFILLER_37_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1165_ clk_divider.count_out\[25\] _0520_ vssd1 vssd1 vccd1 vccd1 _0526_ sky130_fd_sc_hd__or2_1
XFILLER_25_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1096_ _0464_ _0467_ _0468_ net100 vssd1 vssd1 vccd1 vccd1 clk_divider.next_count\[13\]
+ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_82_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_72_Left_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_20_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1376__A net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0949_ _0304_ _0302_ vssd1 vssd1 vccd1 vccd1 _0339_ sky130_fd_sc_hd__and2b_1
XFILLER_69_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_81_Left_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_75_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_47_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_83_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_55_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_54_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_90_Left_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_34_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_50_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_39_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_78_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_66_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_6_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_19_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_62_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_61_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_91_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_30_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0803_ _0170_ _0192_ vssd1 vssd1 vccd1 vccd1 _0193_ sky130_fd_sc_hd__nand2_2
X_0734_ net124 _0123_ vssd1 vssd1 vccd1 vccd1 _0124_ sky130_fd_sc_hd__nand2_1
X_0665_ _0048_ _0054_ vssd1 vssd1 vccd1 vccd1 _0055_ sky130_fd_sc_hd__xnor2_2
XFILLER_97_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_69_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_97_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_68_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1217_ _0350_ _0492_ clk_divider.next_count\[20\] _0330_ _0574_ vssd1 vssd1 vccd1
+ vccd1 _0575_ sky130_fd_sc_hd__a221o_1
XFILLER_65_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_52_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1148_ clk_divider.count_out\[22\] net109 vssd1 vssd1 vccd1 vccd1 _0512_ sky130_fd_sc_hd__or2_1
XFILLER_80_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1079_ clk_divider.count_out\[11\] net93 net91 vssd1 vssd1 vccd1 vccd1 _0454_ sky130_fd_sc_hd__and3_1
XFILLER_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_21_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_91_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_44_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_100_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_101_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_12_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_8_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_61_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_94_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_79_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_39_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_94_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_79_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_94_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_65_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1002_ _0354_ _0391_ _0352_ vssd1 vssd1 vccd1 vccd1 _0392_ sky130_fd_sc_hd__a21o_1
XFILLER_34_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_62_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_77_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0717_ net14 _0086_ vssd1 vssd1 vccd1 vccd1 _0107_ sky130_fd_sc_hd__xnor2_2
XFILLER_89_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0648_ net17 net16 vssd1 vssd1 vccd1 vccd1 _0038_ sky130_fd_sc_hd__xor2_2
XFILLER_97_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_85_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1154__B1 net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_88_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_283 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_13_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_53_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_21_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_5_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput22 net22 vssd1 vssd1 vccd1 vccd1 gpio_oeb[0] sky130_fd_sc_hd__buf_2
Xoutput33 net33 vssd1 vssd1 vccd1 vccd1 gpio_oeb[1] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_8_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput55 net55 vssd1 vssd1 vccd1 vccd1 gpio_oeb[9] sky130_fd_sc_hd__buf_2
Xoutput66 net66 vssd1 vssd1 vccd1 vccd1 gpio_out[19] sky130_fd_sc_hd__buf_2
Xoutput44 net44 vssd1 vssd1 vccd1 vccd1 gpio_oeb[2] sky130_fd_sc_hd__buf_2
XFILLER_88_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
Xoutput77 net77 vssd1 vssd1 vccd1 vccd1 gpio_out[29] sky130_fd_sc_hd__buf_2
Xoutput88 net88 vssd1 vssd1 vccd1 vccd1 gpio_out[8] sky130_fd_sc_hd__buf_2
XFILLER_0_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_76_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_0_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_76_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_29_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_91_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_44_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_62 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_16_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_31_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_70_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_31_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_42_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_99_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_86_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_79_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_67_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_23_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_35_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_50_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_50_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_10_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_50_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_89_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_89_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_58_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_58_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_93_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_45_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_58_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_73_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_26_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_41_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_11_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_1_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_3_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_1_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_49_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_19_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_17_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_32_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_32_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0982_ _0010_ clk_divider.count_out\[7\] vssd1 vssd1 vccd1 vccd1 _0372_ sky130_fd_sc_hd__nand2_1
XFILLER_32_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1054__C1 _0036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_74_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout108 count\[0\] vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__clkbuf_2
Xfanout119 net120 vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__clkbuf_4
XFILLER_101_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xteam_00_129 vssd1 vssd1 vccd1 vccd1 team_00_129/HI la_data_out[3] sky130_fd_sc_hd__conb_1
XFILLER_27_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_82_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_55_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_85_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_70_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_23_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_96_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1318__CLK clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_85_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_73_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_54_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_61_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_14_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_14_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_TAPCELL_ROW_99_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_68_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1250_ _0000_ net105 net108 count\[1\] vssd1 vssd1 vccd1 vccd1 _0598_ sky130_fd_sc_hd__or4b_1
X_1181_ _0537_ _0538_ vssd1 vssd1 vccd1 vccd1 _0539_ sky130_fd_sc_hd__nand2_1
XFILLER_76_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_24_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_37_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_17_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_52_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0965_ _0018_ _0180_ vssd1 vssd1 vccd1 vccd1 _0355_ sky130_fd_sc_hd__xnor2_1
X_0896_ _0250_ _0253_ _0284_ _0285_ vssd1 vssd1 vccd1 vccd1 _0286_ sky130_fd_sc_hd__a211o_1
XFILLER_59_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_74_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_74_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1379_ net115 vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__clkbuf_1
XFILLER_36_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_43_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_55_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_90_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_51_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_21_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__0741__A net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1290__CLK clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_100_Left_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_57_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_64_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_64_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_14_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_9_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_80_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout90 _0403_ vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__buf_2
X_0750_ _0011_ _0012_ _0139_ _0138_ vssd1 vssd1 vccd1 vccd1 _0140_ sky130_fd_sc_hd__o31a_1
XANTENNA__0651__A net18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0681_ net15 _0070_ vssd1 vssd1 vccd1 vccd1 _0071_ sky130_fd_sc_hd__xnor2_1
XFILLER_89_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_71_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1302_ clknet_2_1__leaf_clk clk_divider.next_count\[18\] net120 vssd1 vssd1 vccd1
+ vccd1 clk_divider.count_out\[18\] sky130_fd_sc_hd__dfrtp_1
X_1233_ _0585_ _0587_ vssd1 vssd1 vccd1 vccd1 _0588_ sky130_fd_sc_hd__nor2_1
XFILLER_29_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_96_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_64_120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1164_ clk_divider.count_out\[25\] _0520_ vssd1 vssd1 vccd1 vccd1 _0525_ sky130_fd_sc_hd__nand2_1
XFILLER_92_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_18_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_37_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1095_ clk_divider.count_out\[13\] net111 vssd1 vssd1 vccd1 vccd1 _0468_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_82_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_20_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_20_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0948_ _0016_ _0337_ _0308_ clk_divider.count_out\[25\] vssd1 vssd1 vccd1 vccd1 _0338_
+ sky130_fd_sc_hd__a2bb2o_1
X_0879_ net125 _0003_ vssd1 vssd1 vccd1 vccd1 _0269_ sky130_fd_sc_hd__or2_1
XFILLER_87_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_28_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__0829__A2 net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_55_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__0736__A net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_54_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__1288__RESET_B net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_34_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_50_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_59_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_93_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_78_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_6_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_19_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0646__A net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_61_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0802_ _0165_ _0169_ vssd1 vssd1 vccd1 vccd1 _0192_ sky130_fd_sc_hd__or2_1
XFILLER_30_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0733_ _0120_ _0121_ vssd1 vssd1 vccd1 vccd1 _0123_ sky130_fd_sc_hd__xor2_2
X_0664_ _0042_ _0052_ vssd1 vssd1 vccd1 vccd1 _0054_ sky130_fd_sc_hd__xor2_2
XFILLER_69_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_68_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1216_ _0368_ clk_divider.next_count\[8\] clk_divider.next_count\[19\] _0347_ vssd1
+ vssd1 vccd1 vccd1 _0574_ sky130_fd_sc_hd__o22ai_1
XFILLER_65_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_1_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_52_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1147_ net96 _0509_ _0510_ _0036_ vssd1 vssd1 vccd1 vccd1 _0511_ sky130_fd_sc_hd__a31o_1
XFILLER_80_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_25_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1078_ _0449_ _0452_ _0453_ net101 vssd1 vssd1 vccd1 vccd1 clk_divider.next_count\[10\]
+ sky130_fd_sc_hd__o211a_1
XFILLER_40_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1310__RESET_B net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_88_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_56_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_28_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_61_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_61_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_98_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_226 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_39_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_94_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_65_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1001_ _0018_ _0180_ _0353_ vssd1 vssd1 vccd1 vccd1 _0391_ sky130_fd_sc_hd__or3b_1
XFILLER_62_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_22_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_34_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_77_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0716_ net13 _0105_ _0104_ vssd1 vssd1 vccd1 vccd1 _0106_ sky130_fd_sc_hd__a21boi_2
XFILLER_7_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_0647_ _0007_ _0008_ vssd1 vssd1 vccd1 vccd1 _0037_ sky130_fd_sc_hd__nor2_1
XFILLER_97_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_57_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_88_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_0_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_13_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_80_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_40_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_5_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_8_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput34 net34 vssd1 vssd1 vccd1 vccd1 gpio_oeb[20] sky130_fd_sc_hd__buf_2
Xoutput23 net23 vssd1 vssd1 vccd1 vccd1 gpio_oeb[10] sky130_fd_sc_hd__buf_2
Xoutput45 net45 vssd1 vssd1 vccd1 vccd1 gpio_oeb[30] sky130_fd_sc_hd__buf_2
Xoutput67 net67 vssd1 vssd1 vccd1 vccd1 gpio_out[1] sky130_fd_sc_hd__buf_2
Xoutput56 net56 vssd1 vssd1 vccd1 vccd1 gpio_out[0] sky130_fd_sc_hd__buf_2
Xoutput89 net89 vssd1 vssd1 vccd1 vccd1 gpio_out[9] sky130_fd_sc_hd__buf_2
Xoutput78 net78 vssd1 vssd1 vccd1 vccd1 gpio_out[2] sky130_fd_sc_hd__buf_2
XFILLER_76_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_76_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_91_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA_input16_A prescaler[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_44_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_56_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_71_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_clkbuf_2_0__f_clk_X clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_72_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_72_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_8_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_98_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_97_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_79_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_94_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_67_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_39_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_94_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_47_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_62_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_50_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_22_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_89_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_77_19 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA_input8_A prescaler[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_97_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_58_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_73_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_26_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_14_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_11_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_42_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_1_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_3_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_76_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_1_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_49_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_91_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input19_X net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_47_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_32_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_44_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0981_ clk_divider.count_out\[8\] _0368_ vssd1 vssd1 vccd1 vccd1 _0371_ sky130_fd_sc_hd__nor2_1
XFILLER_8_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_59_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_74_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout109 net110 vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__buf_2
XFILLER_79_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_94_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_85_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_50_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_96_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_58_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_58_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_100_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_24_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_40 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_1_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_68_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1180_ _0193_ clk_divider.next_count\[10\] vssd1 vssd1 vccd1 vccd1 _0538_ sky130_fd_sc_hd__xor2_1
XFILLER_37_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_94_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_91_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_32_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_32_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_60_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0964_ clk_divider.count_out\[17\] _0179_ vssd1 vssd1 vccd1 vccd1 _0354_ sky130_fd_sc_hd__nand2_1
X_0895_ _0233_ _0266_ vssd1 vssd1 vccd1 vccd1 _0285_ sky130_fd_sc_hd__or2_1
XFILLER_99_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_101_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_87_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_4_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1378_ net116 vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__clkbuf_1
XFILLER_83_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_195 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_55_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_11_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_51_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_11_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_23_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_21_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_48_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_29_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_57_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_61_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_14_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_9_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_42_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout91 _0403_ vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__clkbuf_2
XFILLER_80_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__0651__B net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0680_ _0058_ _0068_ vssd1 vssd1 vccd1 vccd1 _0070_ sky130_fd_sc_hd__xor2_1
XFILLER_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_69_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1301_ clknet_2_0__leaf_clk clk_divider.next_count\[17\] net120 vssd1 vssd1 vccd1
+ vccd1 clk_divider.count_out\[17\] sky130_fd_sc_hd__dfrtp_1
XFILLER_84_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1232_ count\[5\] net107 _0579_ _0586_ vssd1 vssd1 vccd1 vccd1 _0587_ sky130_fd_sc_hd__o31ai_2
XFILLER_64_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1163_ clk_divider.count_out\[25\] net92 net90 vssd1 vssd1 vccd1 vccd1 _0524_ sky130_fd_sc_hd__and3_1
XFILLER_64_176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_52_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1094_ net94 _0465_ _0466_ net111 vssd1 vssd1 vccd1 vccd1 _0467_ sky130_fd_sc_hd__o31ai_1
XTAP_TAPCELL_ROW_82_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_100_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_33_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1308__CLK clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0947_ _0015_ _0298_ _0307_ _0311_ vssd1 vssd1 vccd1 vccd1 _0337_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout116_A net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0878_ net11 net125 vssd1 vssd1 vccd1 vccd1 _0268_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_93_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_28_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_83_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_26_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_54_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_34_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xclkload0 clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload0/X sky130_fd_sc_hd__clkbuf_4
XFILLER_50_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_3_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_75 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_66_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_6_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_75_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_34_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0646__B net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_61_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_91_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_15_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_30_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0801_ _0171_ _0190_ vssd1 vssd1 vccd1 vccd1 _0191_ sky130_fd_sc_hd__or2_2
X_0732_ _0120_ _0121_ vssd1 vssd1 vccd1 vccd1 _0122_ sky130_fd_sc_hd__nand2_1
X_0663_ _0042_ _0052_ vssd1 vssd1 vccd1 vccd1 _0053_ sky130_fd_sc_hd__nor2_1
XFILLER_41_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_69_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1215_ _0179_ clk_divider.next_count\[17\] _0571_ _0572_ vssd1 vssd1 vccd1 vccd1
+ _0573_ sky130_fd_sc_hd__o211ai_1
XFILLER_25_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_37_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1146_ clk_divider.count_out\[22\] _0503_ vssd1 vssd1 vccd1 vccd1 _0510_ sky130_fd_sc_hd__or2_1
XFILLER_80_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_65_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_1_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_25_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_80_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1077_ clk_divider.count_out\[10\] net112 vssd1 vssd1 vccd1 vccd1 _0453_ sky130_fd_sc_hd__or2_1
XFILLER_33_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_31_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_96_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_88_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_0_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_16_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_39_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_43_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_94_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_66_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_47_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_59_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_81_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1000_ _0349_ _0350_ clk_divider.count_out\[18\] vssd1 vssd1 vccd1 vccd1 _0390_ sky130_fd_sc_hd__or3b_1
XFILLER_19_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_47_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_62_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_50_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_89_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_30_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_0_clk_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0715_ _0102_ _0103_ vssd1 vssd1 vccd1 vccd1 _0105_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_77_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0646_ net118 net4 net2 vssd1 vssd1 vccd1 vccd1 _0036_ sky130_fd_sc_hd__or3b_4
XFILLER_97_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_85_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_69_Left_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_65_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_36_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1129_ net96 _0494_ _0495_ _0036_ vssd1 vssd1 vccd1 vccd1 _0496_ sky130_fd_sc_hd__a31o_1
XFILLER_15_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_21_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_EDGE_ROW_78_Left_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_31_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
Xoutput24 net24 vssd1 vssd1 vccd1 vccd1 gpio_oeb[11] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_8_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput46 net46 vssd1 vssd1 vccd1 vccd1 gpio_oeb[31] sky130_fd_sc_hd__buf_2
Xoutput57 net57 vssd1 vssd1 vccd1 vccd1 gpio_out[10] sky130_fd_sc_hd__buf_2
Xoutput35 net35 vssd1 vssd1 vccd1 vccd1 gpio_oeb[21] sky130_fd_sc_hd__buf_2
Xoutput79 net79 vssd1 vssd1 vccd1 vccd1 gpio_out[30] sky130_fd_sc_hd__buf_2
XFILLER_0_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput68 net68 vssd1 vssd1 vccd1 vccd1 gpio_out[20] sky130_fd_sc_hd__buf_2
XFILLER_88_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_76_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_91_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_29_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_29_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_19_Right_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_31_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_44_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_31_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_70_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_42_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_8_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_99_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_EDGE_ROW_28_Right_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_67_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_94_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_39_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_94_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_37_Right_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_50_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_30_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_46_Right_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_89_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_89_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0629_ net106 net107 vssd1 vssd1 vccd1 vccd1 _0022_ sky130_fd_sc_hd__and2_1
XFILLER_58_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_97_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_85_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_55_Right_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_26_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_81_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_26_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_13_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_41_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_64_Right_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0760__A net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_5_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_3_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_49_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_73_Right_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__0638__C clk_divider.rollover_flag vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_82_Right_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0980_ _0369_ vssd1 vssd1 vccd1 vccd1 _0370_ sky130_fd_sc_hd__inv_2
XFILLER_32_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_12_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_8_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_74_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_101_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_91_Right_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_300 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_94_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_55_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_85_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_23_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_12_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_96_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout101_X net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_58_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_44_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_24_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_52_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_96_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_78_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_1_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_49_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_91_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_45_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_60_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_20_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0963_ clk_divider.count_out\[17\] _0179_ vssd1 vssd1 vccd1 vccd1 _0353_ sky130_fd_sc_hd__or2_1
XFILLER_9_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0894_ _0279_ _0283_ vssd1 vssd1 vccd1 vccd1 _0284_ sky130_fd_sc_hd__or2_1
XFILLER_99_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_101_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1377_ net115 vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__clkbuf_1
XFILLER_95_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1304__RESET_B net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_11_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_23_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_98_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_21_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_74_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_19_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_48_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_100_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_29_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_61_306 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_64_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_14_Left_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_9_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_14_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_80_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout92 net95 vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__buf_2
XFILLER_6_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_89_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_EDGE_ROW_23_Left_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_71_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1300_ clknet_2_0__leaf_clk clk_divider.next_count\[16\] net119 vssd1 vssd1 vccd1
+ vccd1 clk_divider.count_out\[16\] sky130_fd_sc_hd__dfrtp_2
X_1231_ net1 _0024_ _0025_ vssd1 vssd1 vccd1 vccd1 _0586_ sky130_fd_sc_hd__and3_1
XFILLER_1_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_77_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1162_ _0519_ _0522_ _0523_ net98 vssd1 vssd1 vccd1 vccd1 clk_divider.next_count\[24\]
+ sky130_fd_sc_hd__o211a_1
XFILLER_92_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_32_Left_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1093_ clk_divider.count_out\[12\] _0455_ clk_divider.count_out\[13\] vssd1 vssd1
+ vccd1 vccd1 _0466_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_82_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_45_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_60_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0946_ _0334_ _0335_ _0309_ _0313_ vssd1 vssd1 vccd1 vccd1 _0336_ sky130_fd_sc_hd__a211o_1
XFILLER_9_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_41_Left_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0877_ net125 _0003_ vssd1 vssd1 vccd1 vccd1 _0267_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_93_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_50_Left_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_55_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_54_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_70_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_11_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_34_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload1 clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload1/Y sky130_fd_sc_hd__bufinv_16
XFILLER_1_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_78_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1297__RESET_B net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_87 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_93_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_6_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_75_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_74_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_61_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_15_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_30_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_42_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0800_ _0164_ _0170_ vssd1 vssd1 vccd1 vccd1 _0190_ sky130_fd_sc_hd__and2_1
XFILLER_30_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0731_ _0091_ _0101_ vssd1 vssd1 vccd1 vccd1 _0121_ sky130_fd_sc_hd__xnor2_2
XFILLER_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0662_ net10 _0050_ vssd1 vssd1 vccd1 vccd1 _0052_ sky130_fd_sc_hd__xnor2_2
XFILLER_97_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1166__B1 _0036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_38_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1214_ _0296_ _0310_ clk_divider.next_count\[24\] vssd1 vssd1 vccd1 vccd1 _0572_
+ sky130_fd_sc_hd__or3_1
XFILLER_80_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_53_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1145_ clk_divider.count_out\[22\] _0503_ vssd1 vssd1 vccd1 vccd1 _0509_ sky130_fd_sc_hd__nand2_1
XFILLER_65_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_25_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_52_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1076_ net93 _0450_ _0451_ net112 vssd1 vssd1 vccd1 vccd1 _0452_ sky130_fd_sc_hd__o31ai_1
XFILLER_80_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_21_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_40_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_21_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_TAPCELL_ROW_31_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0929_ _0316_ _0317_ clk_divider.count_out\[23\] vssd1 vssd1 vccd1 vccd1 _0319_ sky130_fd_sc_hd__a21oi_1
XFILLER_88_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_88_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_29_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_90_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_67_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_39_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_28_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_43_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_71_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_24_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_100_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_79_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_66_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_86_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_35_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_62_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_62_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_15_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_22_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0714_ _0102_ _0103_ vssd1 vssd1 vccd1 vccd1 _0104_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_77_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0645_ net4 net2 net1 vssd1 vssd1 vccd1 vccd1 _0035_ sky130_fd_sc_hd__and3b_2
XTAP_TAPCELL_ROW_90_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_TAPCELL_ROW_0_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1128_ clk_divider.count_out\[19\] _0488_ vssd1 vssd1 vccd1 vccd1 _0495_ sky130_fd_sc_hd__or2_1
XFILLER_25_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_36_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1059_ clk_divider.count_out\[7\] _0431_ vssd1 vssd1 vccd1 vccd1 _0438_ sky130_fd_sc_hd__or2_1
XFILLER_15_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_25_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
Xoutput25 net25 vssd1 vssd1 vccd1 vccd1 gpio_oeb[12] sky130_fd_sc_hd__buf_2
Xoutput47 net47 vssd1 vssd1 vccd1 vccd1 gpio_oeb[32] sky130_fd_sc_hd__buf_2
Xoutput36 net36 vssd1 vssd1 vccd1 vccd1 gpio_oeb[22] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_8_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput58 net58 vssd1 vssd1 vccd1 vccd1 gpio_out[11] sky130_fd_sc_hd__buf_2
Xoutput69 net69 vssd1 vssd1 vccd1 vccd1 gpio_out[21] sky130_fd_sc_hd__buf_2
XANTENNA__0758__A net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_84_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_17_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_44_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_56_88 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_44_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_44_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_70_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_4_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_94_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_67_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_94_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_6_Left_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_82_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_35_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0628_ count\[4\] net103 net104 count\[5\] vssd1 vssd1 vccd1 vccd1 _0021_ sky130_fd_sc_hd__or4b_1
XFILLER_100_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_97_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_85_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_66_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_26_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_26_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_81_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_26_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_21_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_5_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_5_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_101_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_95_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1293__CLK clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_76_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_49_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_64_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_19_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_36_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_47_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_17_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_9_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__0670__B net18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_74_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_97_Left_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_67_312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_94_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_67_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_55_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_94_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_85_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_10_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_50_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_2_1__f_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_58_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_100_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_37_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_46_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_73_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_26_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_44_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_78 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_24_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_78_64 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_77_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_94_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_92_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_37_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_49_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_91_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_32_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__0681__A net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0962_ _0351_ _0349_ _0348_ vssd1 vssd1 vccd1 vccd1 _0352_ sky130_fd_sc_hd__or3b_1
XFILLER_32_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_60_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_9_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0893_ _0281_ _0282_ vssd1 vssd1 vccd1 vccd1 _0283_ sky130_fd_sc_hd__nand2_1
XFILLER_99_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1376_ net117 vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__clkbuf_1
XFILLER_67_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_83_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_112 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_55_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_23_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_98_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_86_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_58_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_29_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_27_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_14_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_14_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_9_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_42_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout93 net94 vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__buf_2
XFILLER_13_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_10_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_6_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_71_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1230_ _0582_ count\[5\] net1 _0584_ vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__and4bb_1
XFILLER_1_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_49_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_65_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1161_ clk_divider.count_out\[24\] net109 vssd1 vssd1 vccd1 vccd1 _0523_ sky130_fd_sc_hd__or2_1
XFILLER_92_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_37_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_52_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1092_ clk_divider.count_out\[13\] clk_divider.count_out\[12\] _0455_ vssd1 vssd1
+ vccd1 vccd1 _0465_ sky130_fd_sc_hd__and3_1
XFILLER_18_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_82_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0945_ _0319_ _0322_ _0320_ vssd1 vssd1 vccd1 vccd1 _0335_ sky130_fd_sc_hd__o21ba_1
X_0876_ _0264_ _0265_ vssd1 vssd1 vccd1 vccd1 _0266_ sky130_fd_sc_hd__or2_1
XFILLER_9_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_93_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_68_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_95_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1359_ net114 vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__clkbuf_1
XFILLER_55_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_54_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_11_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_34_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload2 clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload2/Y sky130_fd_sc_hd__clkinv_2
XFILLER_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_6_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_75_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_19_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_34_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_30_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0730_ _0010_ _0011_ _0119_ _0118_ vssd1 vssd1 vccd1 vccd1 _0120_ sky130_fd_sc_hd__o31ai_2
X_0661_ net10 _0050_ vssd1 vssd1 vccd1 vccd1 _0051_ sky130_fd_sc_hd__nand2_1
XFILLER_97_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1213_ _0183_ _0476_ clk_divider.next_count\[27\] _0299_ vssd1 vssd1 vccd1 vccd1
+ _0571_ sky130_fd_sc_hd__o22a_1
XFILLER_27_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_38_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_77_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_38_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1144_ clk_divider.count_out\[22\] net92 net90 vssd1 vssd1 vccd1 vccd1 _0508_ sky130_fd_sc_hd__and3_1
XFILLER_80_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1075_ clk_divider.count_out\[9\] _0443_ clk_divider.count_out\[10\] vssd1 vssd1
+ vccd1 vccd1 _0451_ sky130_fd_sc_hd__a21oi_1
XFILLER_25_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_80_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_33_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_21_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout121_A net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0928_ _0316_ _0317_ vssd1 vssd1 vccd1 vccd1 _0318_ sky130_fd_sc_hd__nand2_1
X_0859_ _0088_ _0177_ vssd1 vssd1 vccd1 vccd1 _0249_ sky130_fd_sc_hd__and2b_1
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_88_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_75_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_29_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_29_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_67_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_43_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_45_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_101_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_101_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_100_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_6_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_3_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_86_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_59_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_74_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_34_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_30_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_30_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0713_ _0073_ _0082_ vssd1 vssd1 vccd1 vccd1 _0103_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_77_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0644_ _0001_ _0024_ _0028_ _0034_ vssd1 vssd1 vccd1 vccd1 counter_to_35.next_count\[5\]
+ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_90_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_38_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1127_ clk_divider.count_out\[19\] _0488_ vssd1 vssd1 vccd1 vccd1 _0494_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_64_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1058_ clk_divider.count_out\[7\] _0431_ vssd1 vssd1 vccd1 vccd1 _0437_ sky130_fd_sc_hd__nand2_1
XFILLER_15_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_33_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_31_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_8_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_1_Right_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput37 net37 vssd1 vssd1 vccd1 vccd1 gpio_oeb[23] sky130_fd_sc_hd__buf_2
Xoutput48 net114 vssd1 vssd1 vccd1 vccd1 gpio_oeb[33] sky130_fd_sc_hd__buf_2
Xoutput26 net26 vssd1 vssd1 vccd1 vccd1 gpio_oeb[13] sky130_fd_sc_hd__buf_2
XFILLER_88_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
Xoutput59 net59 vssd1 vssd1 vccd1 vccd1 gpio_out[12] sky130_fd_sc_hd__buf_2
XFILLER_0_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_88_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_48_229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_56_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_56_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_71_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_72_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_4_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_67_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_94_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_47_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_62_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_90_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_15_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_13_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0627_ clk_divider.count_out\[5\] vssd1 vssd1 vccd1 vccd1 _0020_ sky130_fd_sc_hd__inv_2
XFILLER_100_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_85_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_26_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_38_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_26_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_41_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_53_243 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_81_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_41_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_5_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_1_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_67_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_91_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_29_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_input14_A prescaler[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_44_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_47_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_72_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_10_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_99_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_74_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_67_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_94_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_94_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_82_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_85_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_23_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_63_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_23_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_96_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA_input6_A nrst vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_58_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_85_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_26_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_37_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_44_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_54_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_5_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_96_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_91_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA_input17_X net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_45_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_45_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_60_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0961_ clk_divider.count_out\[18\] _0350_ vssd1 vssd1 vccd1 vccd1 _0351_ sky130_fd_sc_hd__xor2_1
XFILLER_20_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0892_ _0258_ _0261_ _0280_ vssd1 vssd1 vccd1 vccd1 _0282_ sky130_fd_sc_hd__nand3_1
XFILLER_9_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_57_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_99_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1375_ net116 vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__clkbuf_1
XFILLER_67_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_82_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_82_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_82_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_23_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1283__CLK clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1313__RESET_B net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_29_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_27_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_42_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_6_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
Xfanout94 net95 vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__buf_2
XFILLER_13_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_6_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_6_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_96_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_49_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_37_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1160_ net92 _0520_ _0521_ net109 vssd1 vssd1 vccd1 vccd1 _0522_ sky130_fd_sc_hd__o31ai_1
XFILLER_92_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_77_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_37_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_92_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1091_ clk_divider.count_out\[13\] net94 net90 vssd1 vssd1 vccd1 vccd1 _0464_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_82_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_60_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_20_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0944_ _0319_ _0320_ _0323_ _0333_ vssd1 vssd1 vccd1 vccd1 _0334_ sky130_fd_sc_hd__or4_1
X_0875_ _0227_ _0229_ _0263_ vssd1 vssd1 vccd1 vccd1 _0265_ sky130_fd_sc_hd__nor3b_1
XTAP_TAPCELL_ROW_93_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_87_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_28_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1358_ net118 vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__clkbuf_1
XFILLER_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1289_ clknet_2_1__leaf_clk clk_divider.next_count\[5\] net120 vssd1 vssd1 vccd1
+ vccd1 clk_divider.count_out\[5\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_26_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_34_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_11_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_34_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_11_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_78_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_6_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_59_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_74_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_59_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_19_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_74_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_62_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_42_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_clkbuf_2_3__f_clk_X clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_6_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0660_ net19 net18 vssd1 vssd1 vccd1 vccd1 _0050_ sky130_fd_sc_hd__xor2_2
XFILLER_97_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1212_ _0013_ clk_divider.next_count\[4\] _0567_ _0568_ _0569_ vssd1 vssd1 vccd1
+ vccd1 _0570_ sky130_fd_sc_hd__o2111ai_1
XFILLER_77_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_77_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1143_ _0507_ vssd1 vssd1 vccd1 vccd1 clk_divider.next_count\[21\] sky130_fd_sc_hd__inv_2
X_1074_ clk_divider.count_out\[10\] clk_divider.count_out\[9\] _0443_ vssd1 vssd1
+ vccd1 vccd1 _0450_ sky130_fd_sc_hd__and3_1
XFILLER_53_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_80_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_21_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_60_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_31_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0927_ _0281_ _0315_ _0279_ vssd1 vssd1 vccd1 vccd1 _0317_ sky130_fd_sc_hd__a21bo_1
X_0858_ _0241_ _0247_ vssd1 vssd1 vccd1 vccd1 _0248_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout114_A net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0789_ _0089_ _0178_ vssd1 vssd1 vccd1 vccd1 _0179_ sky130_fd_sc_hd__xnor2_2
XFILLER_88_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_88_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_67_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_43_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_56_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_71_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_45_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_24_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_101_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_12_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_61_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_8_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_66_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_59_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_74_274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_35_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_62_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_15_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_30_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_42_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_51_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0712_ _0009_ _0010_ _0101_ _0100_ vssd1 vssd1 vccd1 vccd1 _0102_ sky130_fd_sc_hd__o31ai_2
XTAP_TAPCELL_ROW_77_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0643_ clk_divider.rollover_flag _0022_ _0033_ count\[5\] vssd1 vssd1 vccd1 vccd1
+ _0034_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_90_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_29_Left_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_38_400 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_38_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1025__B net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1126_ clk_divider.count_out\[19\] net95 net90 vssd1 vssd1 vccd1 vccd1 _0493_ sky130_fd_sc_hd__and3_1
XFILLER_65_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_0_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_38_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_88_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_36_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1057_ clk_divider.count_out\[7\] net94 net91 vssd1 vssd1 vccd1 vccd1 _0436_ sky130_fd_sc_hd__and3_1
XFILLER_15_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_38_Left_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_31_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA_fanout117_X net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput27 net27 vssd1 vssd1 vccd1 vccd1 gpio_oeb[14] sky130_fd_sc_hd__buf_2
Xoutput38 net38 vssd1 vssd1 vccd1 vccd1 gpio_oeb[24] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_8_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput49 net49 vssd1 vssd1 vccd1 vccd1 gpio_oeb[3] sky130_fd_sc_hd__buf_2
XFILLER_88_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_0_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_88_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_71_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_44_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_72_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_24_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_99_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_21_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_79_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_75_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_90_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0684__B net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_50_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_87_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_30_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_13_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_0626_ clk_divider.count_out\[6\] vssd1 vssd1 vccd1 vccd1 _0019_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_15_Right_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_81_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_EDGE_ROW_24_Right_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_53_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1109_ clk_divider.count_out\[16\] _0474_ vssd1 vssd1 vccd1 vccd1 _0479_ sky130_fd_sc_hd__nor2_1
XFILLER_81_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_41_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_53_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_EDGE_ROW_33_Right_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_1_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_91_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_57_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_72_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_42_Right_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_32_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_12_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_73_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_51_Right_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_99_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_74_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_94_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_60_Right_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_18_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_23_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_35_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_96_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0609_ clk_divider.count_out\[0\] vssd1 vssd1 vccd1 vccd1 _0002_ sky130_fd_sc_hd__inv_2
XFILLER_86_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_100_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_85_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_73_306 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_39_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_54_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_81_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_14_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_41_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_52_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_89_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_78_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_76_111 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_94_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_91_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_76_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_91_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_27_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_45_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_57_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_60_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_60_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0960_ _0241_ _0345_ vssd1 vssd1 vccd1 vccd1 _0350_ sky130_fd_sc_hd__xnor2_2
XFILLER_13_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_60_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_80_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0891_ _0258_ _0261_ _0280_ vssd1 vssd1 vccd1 vccd1 _0281_ sky130_fd_sc_hd__a21o_1
XFILLER_99_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_4_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_68_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_4_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1374_ net117 vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__clkbuf_1
XFILLER_67_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_55_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_82_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_70_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_36_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_51_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_98_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_21_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_64_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1111__B1 net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_42_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_42_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_80_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xfanout95 _0395_ vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_6_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_77_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_37_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_92_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_18_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1090_ _0463_ vssd1 vssd1 vccd1 vccd1 clk_divider.next_count\[12\] sky130_fd_sc_hd__inv_2
XFILLER_92_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_33_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_52_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_82_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_54_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_0943_ _0328_ _0332_ _0327_ vssd1 vssd1 vccd1 vccd1 _0333_ sky130_fd_sc_hd__o21ba_1
X_0874_ _0227_ _0229_ _0263_ vssd1 vssd1 vccd1 vccd1 _0264_ sky130_fd_sc_hd__o21ba_1
XFILLER_9_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_93_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_10_Left_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1357_ net114 vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__clkbuf_1
XFILLER_95_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_68_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1288_ clknet_2_1__leaf_clk clk_divider.next_count\[4\] net120 vssd1 vssd1 vccd1
+ vccd1 clk_divider.count_out\[4\] sky130_fd_sc_hd__dfrtp_2
XFILLER_24_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_26_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_54_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_24_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_34_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_3_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_3_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_101_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_74_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_6_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_47_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_75_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_74_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_74_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_15_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_34_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_91_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_6_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_40_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_97_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1211_ _0368_ clk_divider.next_count\[8\] vssd1 vssd1 vccd1 vccd1 _0569_ sky130_fd_sc_hd__nand2_1
XFILLER_65_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1142_ _0502_ _0505_ _0506_ vssd1 vssd1 vccd1 vccd1 _0507_ sky130_fd_sc_hd__a21o_1
XFILLER_37_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_92_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1073_ clk_divider.count_out\[10\] net93 net91 vssd1 vssd1 vccd1 vccd1 _0449_ sky130_fd_sc_hd__and3_1
XFILLER_18_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_52_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_21_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0926_ _0279_ _0281_ _0315_ vssd1 vssd1 vccd1 vccd1 _0316_ sky130_fd_sc_hd__nand3b_1
X_0857_ _0243_ _0244_ vssd1 vssd1 vccd1 vccd1 _0247_ sky130_fd_sc_hd__xnor2_2
XFILLER_20_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0788_ _0127_ _0175_ _0177_ _0108_ vssd1 vssd1 vccd1 vccd1 _0178_ sky130_fd_sc_hd__a31o_1
XFILLER_0_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_89_Right_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_96_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_68_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_67_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_16_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_39_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_56_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1078__C1 net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_98_Right_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_20_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__1296__CLK clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_101_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_47_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_19_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_74_286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_35_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_30_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_30_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0711_ _0098_ _0099_ vssd1 vssd1 vccd1 vccd1 _0101_ sky130_fd_sc_hd__xnor2_2
XFILLER_11_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_7_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_77_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0642_ count\[4\] net103 net104 vssd1 vssd1 vccd1 vccd1 _0033_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_90_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_97_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_78_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_38_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_38_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_93_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1125_ _0492_ vssd1 vssd1 vccd1 vccd1 clk_divider.next_count\[18\] sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_0_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_88_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1056_ net100 _0434_ _0435_ vssd1 vssd1 vccd1 vccd1 clk_divider.next_count\[6\] sky130_fd_sc_hd__and3_1
XFILLER_33_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_40_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_16_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0909_ _0003_ _0297_ _0200_ vssd1 vssd1 vccd1 vccd1 _0299_ sky130_fd_sc_hd__a21o_1
Xoutput39 net39 vssd1 vssd1 vccd1 vccd1 gpio_oeb[25] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_8_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput28 net28 vssd1 vssd1 vccd1 vccd1 gpio_oeb[15] sky130_fd_sc_hd__buf_2
XFILLER_88_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_88_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_76_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_56_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_71_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_31_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_12_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_8_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_4_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_98_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_79_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_75_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA_clkload2_A clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1311__CLK clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1290__RESET_B net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_15_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_22_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_30_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_13_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_41_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_89_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0625_ clk_divider.count_out\[16\] vssd1 vssd1 vccd1 vccd1 _0018_ sky130_fd_sc_hd__inv_2
XFILLER_58_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_38_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_49_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1108_ clk_divider.count_out\[16\] clk_divider.count_out\[15\] _0469_ vssd1 vssd1
+ vccd1 vccd1 _0478_ sky130_fd_sc_hd__and3_1
X_1039_ clk_divider.count_out\[4\] _0404_ vssd1 vssd1 vccd1 vccd1 _0421_ sky130_fd_sc_hd__nand2_1
XFILLER_13_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_2_Left_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_88_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_57_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_91_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_44_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_72_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_40_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_10_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_57_Left_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_74_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_82_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_66_Left_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_85_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_50_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_75_Left_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_96_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0608_ net1 vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__inv_2
XFILLER_100_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_98_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_84_Left_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_85_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_73_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_39_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_26_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_81_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_26_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_53_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_54_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_93_Left_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_5_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_78_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_77_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_76_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_91_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
Xclkbuf_2_0__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_2_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_60_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_60_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_13_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_43_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0890_ net123 _0275_ vssd1 vssd1 vccd1 vccd1 _0280_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_80_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_4_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_68_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_4_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_68_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1373_ net115 vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__clkbuf_1
XFILLER_4_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_67_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_63_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_36_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_51_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_3_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_48_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_59_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_100_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_46_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1224__B net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_73_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_TAPCELL_ROW_29_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_81_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_42_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_10_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
Xfanout96 _0394_ vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__buf_2
XFILLER_6_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_89_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_92_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_37_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_38_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_64_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_60_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_33_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_13_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0942_ clk_divider.count_out\[20\] _0330_ vssd1 vssd1 vccd1 vccd1 _0332_ sky130_fd_sc_hd__nand2_1
X_0873_ _0261_ _0262_ vssd1 vssd1 vccd1 vccd1 _0263_ sky130_fd_sc_hd__nand2_1
XFILLER_62_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_93_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1356_ net114 vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__clkbuf_1
XFILLER_95_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_18_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1287_ clknet_2_3__leaf_clk clk_divider.next_count\[3\] net119 vssd1 vssd1 vccd1
+ vccd1 clk_divider.count_out\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_55_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_55_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_TAPCELL_ROW_26_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_24_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_24_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_34_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_59_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_86_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_6_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_74_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_46_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_42_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_54_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_42_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_6_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_97_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1210_ net100 _0434_ _0435_ _0011_ vssd1 vssd1 vccd1 vccd1 _0568_ sky130_fd_sc_hd__a31o_1
X_1141_ clk_divider.count_out\[21\] net110 net99 vssd1 vssd1 vccd1 vccd1 _0506_ sky130_fd_sc_hd__o21ai_1
XFILLER_92_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_37_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_92_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_52_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1072_ clk_divider.count_out\[9\] net111 _0445_ _0448_ net100 vssd1 vssd1 vccd1 vccd1
+ clk_divider.next_count\[9\] sky130_fd_sc_hd__o221a_1
XFILLER_45_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_21_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_60_173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_60_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0925_ _0255_ _0288_ _0283_ net102 vssd1 vssd1 vccd1 vccd1 _0315_ sky130_fd_sc_hd__a211o_1
X_0856_ _0243_ _0244_ vssd1 vssd1 vccd1 vccd1 _0246_ sky130_fd_sc_hd__nand2_1
X_0787_ _0106_ _0107_ vssd1 vssd1 vccd1 vccd1 _0177_ sky130_fd_sc_hd__xor2_2
XFILLER_29_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_56_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_67_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_39_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_71_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_45_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_71_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_24_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_101_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_20_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_79_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_10_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_10_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_19_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_74_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1131__C net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_35_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_0710_ _0098_ _0099_ vssd1 vssd1 vccd1 vccd1 _0100_ sky130_fd_sc_hd__nand2_1
XFILLER_11_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_0641_ net103 net104 vssd1 vssd1 vccd1 vccd1 _0032_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_90_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_93_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1124_ _0487_ _0490_ _0491_ vssd1 vssd1 vccd1 vccd1 _0492_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_0_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_53_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_93_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_88_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1055_ clk_divider.count_out\[6\] net112 vssd1 vssd1 vccd1 vccd1 _0435_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_64_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_16_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0908_ _0273_ _0296_ net125 vssd1 vssd1 vccd1 vccd1 _0298_ sky130_fd_sc_hd__o21ai_1
X_0839_ net18 _0228_ vssd1 vssd1 vccd1 vccd1 _0229_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_8_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput29 net29 vssd1 vssd1 vccd1 vccd1 gpio_oeb[16] sky130_fd_sc_hd__buf_2
XFILLER_0_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_56_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_4_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_4_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_97_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_79_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1126__C net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_35_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_90_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_75_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_35_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_46_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_13_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_41_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0624_ clk_divider.count_out\[21\] vssd1 vssd1 vccd1 vccd1 _0017_ sky130_fd_sc_hd__inv_2
XFILLER_97_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_85_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_38_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_66_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_38_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_49_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_5_Right_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1107_ _0018_ net96 _0402_ vssd1 vssd1 vccd1 vccd1 _0477_ sky130_fd_sc_hd__or3_1
X_1038_ _0021_ counter_to_35.next_count\[0\] counter_to_35.next_count\[1\] vssd1 vssd1
+ vccd1 vccd1 counter_to_35.next_flag sky130_fd_sc_hd__and3b_1
XFILLER_22_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__1286__CLK clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout122_X net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_67_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_67_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_17_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_57_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_83_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_72_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_17_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_32_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_12_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_10_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_48_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_18_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_31_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_96_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0607_ clk_divider.rollover_flag vssd1 vssd1 vccd1 vccd1 _0001_ sky130_fd_sc_hd__inv_2
XFILLER_58_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_85_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_100_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_39_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_39_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_54_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_14_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_53_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_81_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_41_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_52_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1301__CLK clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_49_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_89_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_1_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_91_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_input12_A prescaler[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_57_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_72_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_13_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_32_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_13_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_43_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_80_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA_output80_A net80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_4_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1372_ net114 vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__clkbuf_1
XFILLER_83_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_23_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_51_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_90_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_31_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_2_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_86_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA_input4_A la_oenb[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_100_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_86_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_100_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_57_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_81_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_14_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_80_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_10_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
Xfanout97 _0394_ vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_89_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_65_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input15_X net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_92_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_33_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_60_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0941_ clk_divider.count_out\[20\] _0330_ vssd1 vssd1 vccd1 vccd1 _0331_ sky130_fd_sc_hd__and2_1
XFILLER_60_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_13_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0872_ _0005_ _0260_ vssd1 vssd1 vccd1 vccd1 _0262_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_93_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1355_ net116 vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__clkbuf_1
XFILLER_68_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_68_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_83_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1286_ clknet_2_0__leaf_clk clk_divider.next_count\[2\] net119 vssd1 vssd1 vccd1
+ vccd1 clk_divider.count_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_71_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_70_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_26_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_63_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_34_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_51_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_34_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_59_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA_input7_X net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_6_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_74_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_15_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1251__A _0589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_54_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_42_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_54_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_6_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_79_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_2_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_37_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_38_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1284__RESET_B net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1140_ net92 _0503_ _0504_ net110 vssd1 vssd1 vccd1 vccd1 _0505_ sky130_fd_sc_hd__o31a_1
XFILLER_92_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_65_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_53_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1071_ net97 _0446_ _0447_ _0036_ vssd1 vssd1 vccd1 vccd1 _0448_ sky130_fd_sc_hd__a31o_1
XFILLER_92_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_80_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_21_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_60_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_TAPCELL_ROW_31_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0924_ _0255_ _0288_ net102 vssd1 vssd1 vccd1 vccd1 _0314_ sky130_fd_sc_hd__a21oi_1
X_0855_ _0243_ _0244_ vssd1 vssd1 vccd1 vccd1 _0245_ sky130_fd_sc_hd__nor2_1
X_0786_ _0127_ _0175_ vssd1 vssd1 vccd1 vccd1 _0176_ sky130_fd_sc_hd__nand2_1
XFILLER_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_83_200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_3_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1269_ _0593_ _0605_ vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_39_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_83_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_45_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_24_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_36_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_10_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_3_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1246__A _0589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_10_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_87_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_59_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_47_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_35_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_62_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_42_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0640_ _0028_ _0030_ _0031_ vssd1 vssd1 vccd1 vccd1 counter_to_35.next_count\[1\]
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_90_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_93_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1123_ clk_divider.count_out\[18\] net110 net98 vssd1 vssd1 vccd1 vccd1 _0491_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_0_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_93_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_88_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1054_ clk_divider.count_out\[6\] _0404_ _0433_ net97 _0036_ vssd1 vssd1 vccd1 vccd1
+ _0434_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_64_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_18_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_16_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0907_ _0286_ _0290_ _0295_ vssd1 vssd1 vccd1 vccd1 _0297_ sky130_fd_sc_hd__a21o_1
X_0838_ _0224_ _0226_ vssd1 vssd1 vccd1 vccd1 _0228_ sky130_fd_sc_hd__xnor2_1
X_0769_ _0149_ _0157_ vssd1 vssd1 vccd1 vccd1 _0159_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_8_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_84_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_24_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_40_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_76_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_87_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_90_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_75_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_35_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_47_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_90_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_43_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_30_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_62_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_41_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0623_ clk_divider.count_out\[24\] vssd1 vssd1 vccd1 vccd1 _0016_ sky130_fd_sc_hd__inv_2
XFILLER_98_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_97_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_66_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_93_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_81_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1106_ _0476_ vssd1 vssd1 vccd1 vccd1 clk_divider.next_count\[15\] sky130_fd_sc_hd__inv_2
XFILLER_26_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_49_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1037_ _0028_ _0419_ _0420_ vssd1 vssd1 vccd1 vccd1 counter_to_35.next_count\[4\]
+ sky130_fd_sc_hd__and3_1
XFILLER_22_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1316__RESET_B net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_88_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_76_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_67_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_84_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_17_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_29_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_83_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_72_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_72_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_16_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_25_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_13_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_EDGE_ROW_11_Right_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_12_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_40_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_4_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_20_Right_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_48_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_63_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_46_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_31_475 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_96_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0606_ count\[3\] vssd1 vssd1 vccd1 vccd1 _0000_ sky130_fd_sc_hd__inv_2
XFILLER_98_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_100_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_37_18 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_39_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_85_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1123__B1 net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_39_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_54_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_54_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_41_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_53_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__1254__A _0589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_64_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_45_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_17_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_27_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_13_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_23_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1371_ net118 vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__clkbuf_1
XFILLER_95_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_48_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_75_191 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_23_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_36_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_51_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_86_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_59_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_86_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_58_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_86_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_73_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_46_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_57_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_10_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
Xfanout98 net101 vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__buf_2
XFILLER_50_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_10_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_20_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1249__A _0589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_89_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1299__CLK clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_8_Left_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_1_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_18_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_49_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_64_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1099__C1 _0036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_57_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_82_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_33_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0940_ _0254_ _0329_ vssd1 vssd1 vccd1 vccd1 _0330_ sky130_fd_sc_hd__or2_1
XFILLER_13_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_20_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_60_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_9_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0871_ _0005_ _0260_ vssd1 vssd1 vccd1 vccd1 _0261_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_93_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_68_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_68_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1354_ net114 vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__clkbuf_1
XFILLER_68_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_28_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1285_ clknet_2_3__leaf_clk clk_divider.next_count\[1\] net119 vssd1 vssd1 vccd1
+ vccd1 clk_divider.count_out\[1\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_54_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_34_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_59_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_101_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_75_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_61_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_91_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_24_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_30_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_24_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_10_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_79_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_49_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1314__CLK clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1070_ clk_divider.count_out\[9\] _0443_ vssd1 vssd1 vccd1 vccd1 _0447_ sky130_fd_sc_hd__or2_1
XFILLER_92_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_65_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_33_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_31_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0923_ clk_divider.count_out\[25\] _0308_ _0312_ _0302_ _0305_ vssd1 vssd1 vccd1
+ vccd1 _0313_ sky130_fd_sc_hd__a2111o_1
X_0854_ net17 _0222_ vssd1 vssd1 vccd1 vccd1 _0244_ sky130_fd_sc_hd__xnor2_2
X_0785_ _0147_ _0173_ _0128_ _0146_ vssd1 vssd1 vccd1 vccd1 _0175_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_49_Right_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_68_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_3_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1268_ _0592_ _0605_ vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_39_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_58_Right_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1199_ _0191_ clk_divider.next_count\[11\] vssd1 vssd1 vccd1 vccd1 _0557_ sky130_fd_sc_hd__nor2_1
XFILLER_24_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_43_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_101_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_12_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_51_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_EDGE_ROW_67_Right_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_3_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_79_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_10_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_87_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_98_Left_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_76_Right_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_34_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_35_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_42_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_70_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_85_Right_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_94_Right_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1122_ net95 _0488_ _0489_ net110 vssd1 vssd1 vccd1 vccd1 _0490_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_0_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1053_ _0431_ _0432_ vssd1 vssd1 vccd1 vccd1 _0433_ sky130_fd_sc_hd__nor2_1
XFILLER_65_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_36_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_80_259 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_21_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_61_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_16_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0906_ _0286_ _0290_ _0295_ vssd1 vssd1 vccd1 vccd1 _0296_ sky130_fd_sc_hd__a21oi_2
X_0837_ _0226_ _0224_ vssd1 vssd1 vccd1 vccd1 _0227_ sky130_fd_sc_hd__and2b_1
X_0768_ _0157_ _0149_ vssd1 vssd1 vccd1 vccd1 _0158_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_8_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0699_ _0088_ vssd1 vssd1 vccd1 vccd1 _0089_ sky130_fd_sc_hd__inv_2
XFILLER_69_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_84_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_72_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_24_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_52_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_4_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__1257__A _0589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_97_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_79_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_94_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_35_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_90_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_46_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_13_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_7_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_0622_ clk_divider.count_out\[25\] vssd1 vssd1 vccd1 vccd1 _0015_ sky130_fd_sc_hd__inv_2
XFILLER_98_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_97_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_85_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_38_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_93_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_66_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_49_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1105_ clk_divider.count_out\[15\] net112 _0472_ _0475_ net99 vssd1 vssd1 vccd1 vccd1
+ _0476_ sky130_fd_sc_hd__o221ai_4
XFILLER_81_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1036_ count\[5\] _0001_ _0023_ _0033_ vssd1 vssd1 vccd1 vccd1 _0420_ sky130_fd_sc_hd__or4b_1
XFILLER_34_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__0716__A1 net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_29_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_72_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_17_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_72_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_16_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_17_Left_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_16_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_40_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_12_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_32_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_10_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_4_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_26_Left_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_79_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_79_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_94_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_48_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_18_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_46_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkload0_A clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_63_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_35_Left_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_31_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_78_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_7_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_44_Left_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_96_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_58_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1063__C net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_93_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_53_Left_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1019_ clk_divider.count_out\[0\] clk_divider.count_out\[1\] net111 vssd1 vssd1 vccd1
+ vccd1 _0408_ sky130_fd_sc_hd__and3_1
XFILLER_22_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_6_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_EDGE_ROW_62_Left_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_73_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_76_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_71_Left_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_72_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_17_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_57_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_72_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_45_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_40_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_EDGE_ROW_80_Left_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0614__A net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1370_ net115 vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_36_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_51_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_90_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_98_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_48_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_86_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_100_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_100_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_39_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_39_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_27_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0645__A_N net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xfanout99 net101 vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__buf_2
XFILLER_10_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_6_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_2_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_8_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_65_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_18_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_TAPCELL_ROW_28_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_60_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_72_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_13_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_9_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0870_ _0258_ _0259_ vssd1 vssd1 vccd1 vccd1 _0260_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_93_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_68_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_95_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1353_ net114 vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__clkbuf_1
XFILLER_83_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_68_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1284_ clknet_2_3__leaf_clk clk_divider.next_count\[0\] net121 vssd1 vssd1 vccd1
+ vccd1 clk_divider.count_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_83_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_36_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_54_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0999_ _0352_ _0355_ _0356_ _0388_ vssd1 vssd1 vccd1 vccd1 _0389_ sky130_fd_sc_hd__or4_1
XFILLER_86_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_86_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_101_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_91_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_15_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_25_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_24_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_10_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_24_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_10_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_40_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_79_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_5_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_1_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_18_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_80_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_33_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_14_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1293__RESET_B net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0922_ _0016_ _0311_ vssd1 vssd1 vccd1 vccd1 _0312_ sky130_fd_sc_hd__xnor2_1
X_0853_ net16 _0237_ _0236_ vssd1 vssd1 vccd1 vccd1 _0243_ sky130_fd_sc_hd__a21boi_2
X_0784_ _0147_ _0173_ _0146_ vssd1 vssd1 vccd1 vccd1 _0174_ sky130_fd_sc_hd__a21o_1
XFILLER_68_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_68_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_96_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput1 en vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_67_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1267_ _0590_ _0600_ _0604_ vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_39_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1289__CLK clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1198_ _0012_ clk_divider.next_count\[5\] vssd1 vssd1 vccd1 vccd1 _0556_ sky130_fd_sc_hd__nor2_1
XFILLER_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_101_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_20_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_86_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_87_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_59_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_47_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_74_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_62_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_30_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_11_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_51_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_97_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_90_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_78_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1162__C1 net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1121_ clk_divider.count_out\[18\] _0483_ vssd1 vssd1 vccd1 vccd1 _0489_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_0_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1052_ clk_divider.count_out\[6\] _0427_ vssd1 vssd1 vccd1 vccd1 _0432_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_64_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_21_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_33_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_16_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0905_ _0270_ _0292_ _0294_ vssd1 vssd1 vccd1 vccd1 _0295_ sky130_fd_sc_hd__a21o_1
X_0836_ net10 _0225_ vssd1 vssd1 vccd1 vccd1 _0226_ sky130_fd_sc_hd__xnor2_1
X_0767_ _0155_ _0156_ _0154_ vssd1 vssd1 vccd1 vccd1 _0157_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_8_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_0698_ _0071_ _0087_ vssd1 vssd1 vccd1 vccd1 _0088_ sky130_fd_sc_hd__xnor2_1
XFILLER_69_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_69_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_29_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_84_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_29_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_44_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_12_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_8_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1304__CLK clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_97_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_79_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_101_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_87_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_47_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_87_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_90_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__0617__A net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_15_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_13_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0621_ clk_divider.count_out\[26\] vssd1 vssd1 vccd1 vccd1 _0014_ sky130_fd_sc_hd__inv_2
XFILLER_97_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_23_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_66_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_81_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1104_ net94 _0473_ _0474_ net111 vssd1 vssd1 vccd1 vccd1 _0475_ sky130_fd_sc_hd__o31ai_2
XFILLER_93_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1035_ _0032_ _0415_ count\[4\] vssd1 vssd1 vccd1 vccd1 _0419_ sky130_fd_sc_hd__a21o_1
XFILLER_22_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1358__A net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0819_ _0202_ _0208_ vssd1 vssd1 vccd1 vccd1 _0209_ sky130_fd_sc_hd__nand2_1
XFILLER_1_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_69_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_84_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_72_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_72_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_25_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_44_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_25_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_9_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_40_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_40_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_10_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_32_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_4_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_4_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_79_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_4_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1117__C1 _0036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_63_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_18_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_46_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_35_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_90_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__0643__A1 clk_divider.rollover_flag vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0634__X _0027_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_31_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_96_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_9_Right_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_98_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_85_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_85_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__0809__X _0199_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_93_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_81_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1018_ net111 _0405_ _0406_ _0407_ vssd1 vssd1 vccd1 vccd1 clk_divider.next_count\[0\]
+ sky130_fd_sc_hd__a211oi_1
XFILLER_22_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_22_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA_fanout120_X net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0720__A net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_77_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_94_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_69_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_57_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_84_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_17_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_72_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_25_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_23_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_4_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_68_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_83_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_36_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_84_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_63_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_51_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_90_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_59_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__1371__A net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_27_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_54_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_89_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_20_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_77_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_49_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_38_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_92_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_18_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_38_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_28_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input10_A prescaler[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_33_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_54_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1352_ net116 vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__clkbuf_1
XFILLER_68_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1283_ clknet_2_0__leaf_clk clk_divider.next_flag net119 vssd1 vssd1 vccd1 vccd1
+ clk_divider.rollover_flag sky130_fd_sc_hd__dfrtp_4
XFILLER_95_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_36_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_91_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_36_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_34_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0998_ _0357_ _0359_ _0361_ _0387_ _0358_ vssd1 vssd1 vccd1 vccd1 _0388_ sky130_fd_sc_hd__o221a_1
XFILLER_99_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_101_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_59_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_75_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input2_A la_data_in[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_86_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_74_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_70_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_15_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_54_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_23_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_24_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_10_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_10_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_40_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_79_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_2_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_65_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_5_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input13_X net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_18_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_73_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_18_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0921_ _0296_ _0310_ vssd1 vssd1 vccd1 vccd1 _0311_ sky130_fd_sc_hd__nor2_1
XFILLER_81_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_TAPCELL_ROW_31_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0852_ _0241_ vssd1 vssd1 vccd1 vccd1 _0242_ sky130_fd_sc_hd__inv_2
X_0783_ _0162_ _0172_ _0148_ vssd1 vssd1 vccd1 vccd1 _0173_ sky130_fd_sc_hd__a21oi_2
XFILLER_53_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_5_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_96_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_29_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_68_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
Xinput2 la_data_in[0] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_1
XFILLER_56_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_67_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1266_ _0582_ _0605_ vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_39_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1197_ _0350_ _0492_ _0552_ _0553_ _0554_ vssd1 vssd1 vccd1 vccd1 _0555_ sky130_fd_sc_hd__o2111ai_1
XFILLER_36_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_52_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_101_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_51_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_20_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_59_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_74_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_2_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_42_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_70_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_23_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_7_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1120_ clk_divider.count_out\[18\] _0483_ vssd1 vssd1 vccd1 vccd1 _0488_ sky130_fd_sc_hd__and2_1
XFILLER_65_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1051_ clk_divider.count_out\[6\] _0427_ vssd1 vssd1 vccd1 vccd1 _0431_ sky130_fd_sc_hd__and2_1
XFILLER_65_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_34_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_36_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_61_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_16_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0904_ _0270_ _0293_ _0292_ vssd1 vssd1 vccd1 vccd1 _0294_ sky130_fd_sc_hd__a21oi_1
X_0835_ net123 _0214_ vssd1 vssd1 vccd1 vccd1 _0225_ sky130_fd_sc_hd__nor2_1
X_0766_ _0150_ _0153_ vssd1 vssd1 vccd1 vccd1 _0156_ sky130_fd_sc_hd__xor2_1
X_0697_ net14 _0086_ _0085_ vssd1 vssd1 vccd1 vccd1 _0087_ sky130_fd_sc_hd__a21boi_1
XFILLER_69_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_96_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_69_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_29_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_84_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1318_ clknet_2_2__leaf_clk counter_to_35.next_count\[5\] net122 vssd1 vssd1 vccd1
+ vccd1 count\[5\] sky130_fd_sc_hd__dfrtp_4
XFILLER_84_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1249_ _0589_ _0597_ vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__nor2_1
XFILLER_37_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_72_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_24_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_52_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_76_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1273__B _0605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_87_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_75_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_101_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_62_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_16_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_87_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_62_51 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_13_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_7_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0620_ net7 vssd1 vssd1 vccd1 vccd1 _0013_ sky130_fd_sc_hd__inv_2
XFILLER_97_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_97_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_87_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_78_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_66_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_16_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_66_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_49_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1103_ clk_divider.count_out\[15\] _0469_ vssd1 vssd1 vccd1 vccd1 _0474_ sky130_fd_sc_hd__and2_1
X_1034_ net103 _0416_ _0418_ vssd1 vssd1 vccd1 vccd1 counter_to_35.next_count\[3\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_19_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_81_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_21_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0818_ _0203_ _0207_ vssd1 vssd1 vccd1 vccd1 _0208_ sky130_fd_sc_hd__xnor2_2
XANTENNA_fanout110_A _0035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0749_ _0136_ _0137_ vssd1 vssd1 vccd1 vccd1 _0139_ sky130_fd_sc_hd__xnor2_1
XANTENNA__1374__A net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_69_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_57_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_83_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_40_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_80_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_25_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_40_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1268__B _0605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_40_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1062__C1 net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_79_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_79_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_48_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_94_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_57_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_18_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_46_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_90_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_63_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_73_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_31_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_98_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_100_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_39_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_78_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_81_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1017_ clk_divider.count_out\[0\] net111 net97 vssd1 vssd1 vccd1 vccd1 _0407_ sky130_fd_sc_hd__and3_1
XFILLER_62_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_22_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_22_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__0720__B net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_89_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_17_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_72_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_45_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_32_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_60_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_13_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_40_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_9_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_23_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_4_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1317__CLK clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_59_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_63_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0645__X _0035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_90_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_44_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_83_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_98_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_58_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_14_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_42_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_80_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_22_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_1_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_38_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_38_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_72_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_TAPCELL_ROW_28_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_26_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_33_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_45_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_63 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_79_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1351_ net116 vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__clkbuf_1
XFILLER_95_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1282_ count\[5\] _0579_ _0586_ vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__and3_1
XFILLER_95_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_83_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_36_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_55_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_91_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_24_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_51_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_62_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0997_ _0362_ _0365_ _0366_ _0386_ _0364_ vssd1 vssd1 vccd1 vccd1 _0387_ sky130_fd_sc_hd__o221a_1
XFILLER_99_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1382__A net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_86_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_101_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_86_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_39_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_53_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_82_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_27_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_81_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_59_Left_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_24_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_10_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_10_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_6_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_79_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1276__B _0605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_68_Left_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_77_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_65_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_5_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_18_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_37_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_73_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_18_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_33_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_61_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0920_ _0286_ _0290_ _0295_ vssd1 vssd1 vccd1 vccd1 _0310_ sky130_fd_sc_hd__and3_1
X_0851_ _0238_ _0239_ vssd1 vssd1 vccd1 vccd1 _0241_ sky130_fd_sc_hd__xnor2_2
X_0782_ _0163_ _0171_ vssd1 vssd1 vccd1 vccd1 _0172_ sky130_fd_sc_hd__nand2_1
XFILLER_5_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_46_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_18_Right_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1265_ _0584_ _0587_ vssd1 vssd1 vccd1 vccd1 _0605_ sky130_fd_sc_hd__or2_2
XFILLER_28_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_83_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_67_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput3 la_data_in[1] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_39_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1196_ _0180_ _0482_ vssd1 vssd1 vccd1 vccd1 _0554_ sky130_fd_sc_hd__or2_1
XFILLER_91_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_64_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_101_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_27_Right_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_51_134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_20_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_36_Right_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_2_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_45_Right_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_15_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__0985__A1 net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_54_Right_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_90_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_78_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_93_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1050_ _0426_ _0429_ _0430_ net100 vssd1 vssd1 vccd1 vccd1 clk_divider.next_count\[5\]
+ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_63_Right_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_64_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_34_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_TAPCELL_ROW_36_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_33_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__0813__B net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0903_ net125 _0003_ net11 vssd1 vssd1 vccd1 vccd1 _0293_ sky130_fd_sc_hd__or3b_1
X_0834_ _0212_ _0213_ _0215_ _0218_ vssd1 vssd1 vccd1 vccd1 _0224_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_72_Right_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0765_ net124 _0013_ vssd1 vssd1 vccd1 vccd1 _0155_ sky130_fd_sc_hd__nor2_1
XFILLER_88_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0696_ _0083_ _0084_ vssd1 vssd1 vccd1 vccd1 _0086_ sky130_fd_sc_hd__xor2_2
XFILLER_84_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_81_Right_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1317_ clknet_2_2__leaf_clk counter_to_35.next_count\[4\] net122 vssd1 vssd1 vccd1
+ vccd1 count\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_29_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_84_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1248_ _0000_ _0596_ vssd1 vssd1 vccd1 vccd1 _0597_ sky130_fd_sc_hd__or2_1
XFILLER_71_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1179_ net14 clk_divider.next_count\[7\] vssd1 vssd1 vccd1 vccd1 _0537_ sky130_fd_sc_hd__xnor2_1
XFILLER_52_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_EDGE_ROW_90_Right_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_76_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_7_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_47_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_87_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_41_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_13_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_7_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_3_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_97_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_87_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_66_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_81_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_66_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_49_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1102_ clk_divider.count_out\[15\] _0469_ vssd1 vssd1 vccd1 vccd1 _0473_ sky130_fd_sc_hd__nor2_1
X_1033_ _0032_ _0415_ _0027_ vssd1 vssd1 vccd1 vccd1 _0418_ sky130_fd_sc_hd__a21oi_1
XFILLER_19_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_34_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_21_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1071__B1 _0036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0817_ _0205_ _0206_ vssd1 vssd1 vccd1 vccd1 _0207_ sky130_fd_sc_hd__nor2_1
X_0748_ _0136_ _0137_ vssd1 vssd1 vccd1 vccd1 _0138_ sky130_fd_sc_hd__nand2_1
XFILLER_88_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0679_ _0058_ _0068_ vssd1 vssd1 vccd1 vccd1 _0069_ sky130_fd_sc_hd__nand2_1
XFILLER_84_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_69_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_29_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_57_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_37_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_0_Right_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_12_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_10_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_79_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_48_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_48_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_63_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_18_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_73_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_16_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_43_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_11_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_98_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_98_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_98_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_13_Left_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_39_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_81_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1016_ _0002_ _0036_ _0027_ vssd1 vssd1 vccd1 vccd1 _0406_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_22_Left_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_22_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_31_Left_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_45_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_84_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_EDGE_ROW_40_Left_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_9_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_40_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_23_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_51_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_95_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_4_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_95_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_95_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_67_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_48_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_59_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_84_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_98_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_27_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_66_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_22_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_22_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_50_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_20_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_89_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_77_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_1_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_77_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_92_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1281__C net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_57_151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_28_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_9_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_41_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_70_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_5_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1281_ count\[5\] net107 net1 _0578_ vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__and4_1
XFILLER_95_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_48_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_91_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_36_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_91_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_63_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_51_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_32_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0996_ _0380_ _0384_ _0385_ vssd1 vssd1 vccd1 vccd1 _0386_ sky130_fd_sc_hd__and3_1
XFILLER_99_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_99_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_59_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_101_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_74_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_53_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__0742__A net18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_33_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1307__CLK clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_2_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_6_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_2_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_2_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_49_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_92_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_18_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_73_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_33_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_60_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_33_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_81_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_41_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0850_ _0238_ _0239_ vssd1 vssd1 vccd1 vccd1 _0240_ sky130_fd_sc_hd__nor2_1
X_0781_ _0164_ _0170_ vssd1 vssd1 vccd1 vccd1 _0171_ sky130_fd_sc_hd__nor2_1
XFILLER_5_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_39_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_96_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1264_ _0584_ _0587_ vssd1 vssd1 vccd1 vccd1 _0604_ sky130_fd_sc_hd__nor2_1
XFILLER_56_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_67_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput4 la_oenb[0] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__buf_1
X_1195_ _0421_ _0424_ _0425_ net7 vssd1 vssd1 vccd1 vccd1 _0553_ sky130_fd_sc_hd__a211o_1
XFILLER_36_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_24_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
Xclkbuf_2_1__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_2_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_91_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_51_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_20_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0979_ clk_divider.count_out\[9\] _0195_ _0368_ clk_divider.count_out\[8\] vssd1
+ vssd1 vccd1 vccd1 _0369_ sky130_fd_sc_hd__a22oi_2
XTAP_TAPCELL_ROW_30_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_5_Left_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_99_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_101_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_15_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_27_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_70_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_15_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_23_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_78_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_93_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_18_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_80_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_TAPCELL_ROW_64_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_33_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_92_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0902_ _0201_ _0291_ vssd1 vssd1 vccd1 vccd1 _0292_ sky130_fd_sc_hd__nand2_1
X_0833_ net17 _0222_ vssd1 vssd1 vccd1 vccd1 _0223_ sky130_fd_sc_hd__nand2_1
X_0764_ _0150_ _0153_ vssd1 vssd1 vccd1 vccd1 _0154_ sky130_fd_sc_hd__nor2_1
X_0695_ _0083_ _0084_ vssd1 vssd1 vccd1 vccd1 _0085_ sky130_fd_sc_hd__nand2_1
XFILLER_96_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1316_ clknet_2_2__leaf_clk counter_to_35.next_count\[3\] net122 vssd1 vssd1 vccd1
+ vccd1 count\[3\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_87_Left_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_84_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_2_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1247_ net105 net106 _0580_ net108 vssd1 vssd1 vccd1 vccd1 _0596_ sky130_fd_sc_hd__or4b_1
XFILLER_37_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_37_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1178_ _0184_ clk_divider.next_count\[14\] vssd1 vssd1 vccd1 vccd1 _0536_ sky130_fd_sc_hd__xnor2_1
XFILLER_64_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_52_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_96_Left_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_76_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_7_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_101_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_16_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_87_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_55_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_31_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_13_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_11_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_7_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_3_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_97_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_78_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_93_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_19_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_38_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_49_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1101_ clk_divider.count_out\[15\] net93 net91 vssd1 vssd1 vccd1 vccd1 _0472_ sky130_fd_sc_hd__and3_1
XFILLER_81_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1032_ _0416_ _0417_ vssd1 vssd1 vccd1 vccd1 counter_to_35.next_count\[2\] sky130_fd_sc_hd__nor2_1
XFILLER_19_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_34_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_34_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_21_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_21_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0816_ net11 _0061_ _0204_ vssd1 vssd1 vccd1 vccd1 _0206_ sky130_fd_sc_hd__and3_1
XANTENNA__0840__A net18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0747_ _0114_ _0115_ vssd1 vssd1 vccd1 vccd1 _0137_ sky130_fd_sc_hd__xnor2_1
XFILLER_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_0678_ _0040_ _0067_ vssd1 vssd1 vccd1 vccd1 _0068_ sky130_fd_sc_hd__xor2_1
XFILLER_57_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_29_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_96_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_29_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_84_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_37_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_40_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_10_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1303__RESET_B net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_89_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_87_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_75_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_63_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_73_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_18_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_16_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_31_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0660__A net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_98_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_100_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_66_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_39_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_66_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_19_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1015_ _0002_ net94 net91 _0199_ vssd1 vssd1 vccd1 vccd1 _0405_ sky130_fd_sc_hd__a31o_1
XFILLER_10_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_22_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_89_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_77_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_94_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_57_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_45_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_84_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_40_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_23_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_95_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__0849__A1 net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_48_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_48_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_59_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_90_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1296__RESET_B net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_59_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_98_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_86_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_66_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_27_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_39_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_22_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_50_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_13_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_20_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_89_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_85_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_38_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_28_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_13_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_41_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_9 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_79_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1280_ net107 _0579_ _0587_ vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__nor3_1
XFILLER_0_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_64_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_48_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_91_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_63_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_32_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0995_ clk_divider.count_out\[11\] _0191_ _0381_ vssd1 vssd1 vccd1 vccd1 _0385_ sky130_fd_sc_hd__o21ai_1
XFILLER_99_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_5_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_99_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_59_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_67_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_82_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_50_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_33_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_92_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_49_21 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_77_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_5_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_65_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_1_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_61_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_60_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_41_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0780_ _0165_ _0169_ vssd1 vssd1 vccd1 vccd1 _0170_ sky130_fd_sc_hd__nand2_1
XFILLER_5_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_96_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_96_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_68_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1263_ _0596_ _0601_ vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__nor2_1
Xinput5 la_oenb[1] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__buf_1
XFILLER_49_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_36_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1194_ _0318_ _0518_ vssd1 vssd1 vccd1 vccd1 _0552_ sky130_fd_sc_hd__or2_1
XFILLER_91_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_64_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_101_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_17_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_32_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0978_ _0168_ _0367_ vssd1 vssd1 vccd1 vccd1 _0368_ sky130_fd_sc_hd__nand2_2
XFILLER_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_30_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_99_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_87_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_101_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_19_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_28_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_2_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_15_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_70_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_55_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_30_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_70_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_11_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_7_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_51_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_2_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_78_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_2_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1147__B1 _0036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_78_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_93_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_64_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_46_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_73_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_61_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_14_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0901_ _0003_ _0200_ vssd1 vssd1 vccd1 vccd1 _0291_ sky130_fd_sc_hd__nand2_1
X_0832_ _0211_ _0220_ vssd1 vssd1 vccd1 vccd1 _0222_ sky130_fd_sc_hd__xor2_2
X_0763_ _0008_ _0151_ _0152_ vssd1 vssd1 vccd1 vccd1 _0153_ sky130_fd_sc_hd__or3_1
X_0694_ _0037_ _0057_ vssd1 vssd1 vccd1 vccd1 _0084_ sky130_fd_sc_hd__xnor2_2
XFILLER_51_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_88_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_69_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1315_ clknet_2_2__leaf_clk counter_to_35.next_count\[2\] net122 vssd1 vssd1 vccd1
+ vccd1 count\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_56_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1246_ _0589_ _0595_ vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__nor2_1
XFILLER_25_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1177_ clk_divider.count_out\[27\] net109 _0533_ _0535_ net98 vssd1 vssd1 vccd1 vccd1
+ clk_divider.next_count\[27\] sky130_fd_sc_hd__o221a_1
XFILLER_52_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_92_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_35_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_12_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_52_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_52_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_21_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_76_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1129__B1 _0036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_75_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_87_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_15_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_43_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_2_0__f_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_41_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_87_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_3_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1100_ clk_divider.count_out\[14\] net111 net100 _0471_ vssd1 vssd1 vccd1 vccd1 clk_divider.next_count\[14\]
+ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_49_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1031_ net105 _0415_ _0028_ vssd1 vssd1 vccd1 vccd1 _0417_ sky130_fd_sc_hd__o21ai_1
XFILLER_34_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_74_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_19_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_34_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_99_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_34_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0815_ net11 _0061_ _0204_ vssd1 vssd1 vccd1 vccd1 _0205_ sky130_fd_sc_hd__a21oi_1
X_0746_ _0011_ net124 _0135_ _0133_ vssd1 vssd1 vccd1 vccd1 _0136_ sky130_fd_sc_hd__a31o_1
XFILLER_88_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0677_ _0059_ _0065_ vssd1 vssd1 vccd1 vccd1 _0067_ sky130_fd_sc_hd__xor2_1
XFILLER_84_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_29_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_84_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_57_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_72_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1229_ _0578_ _0583_ vssd1 vssd1 vccd1 vccd1 _0585_ sky130_fd_sc_hd__or2_1
XFILLER_44_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_37_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_25_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_94_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_89_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_57_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input19_A prescaler[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_75_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_18_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_16_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_73_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_16_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_8_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__0660__B net18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_85_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1292__CLK clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_14_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_39_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_81_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_66_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_19_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_54_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1014_ net96 _0402_ vssd1 vssd1 vccd1 vccd1 _0404_ sky130_fd_sc_hd__nor2_2
XFILLER_34_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_8_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0729_ _0116_ _0117_ vssd1 vssd1 vccd1 vccd1 _0119_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_73_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_194 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_69_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_84_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_27_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_38_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_45_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_57_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_84_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_40_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_23_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_51_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_95_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_91_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_75_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_48_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_59_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_36_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_84_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_90_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_16_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_31_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_98_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_66_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_81_123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_81_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_13_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_22_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_22_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_50_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_2_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_77_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_49_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_73_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_56_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_70_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_95_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_95_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_63_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_81_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_32_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0994_ _0369_ _0379_ _0383_ vssd1 vssd1 vccd1 vccd1 _0384_ sky130_fd_sc_hd__a21o_1
XFILLER_5_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_59_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_101_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_19_Left_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_27_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_54_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_28_Left_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_49_33 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_77_259 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_100_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_69_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_5_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_45_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_33_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_60_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__0988__A1 net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_96_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_96_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1262_ _0594_ _0601_ vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__nor2_1
Xinput6 nrst vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__buf_1
XFILLER_76_270 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_37_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_64_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1193_ _0183_ _0476_ clk_divider.next_count\[19\] _0347_ _0550_ vssd1 vssd1 vccd1
+ vccd1 _0551_ sky130_fd_sc_hd__a221o_1
XFILLER_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_36_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_51_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_20_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0977_ net15 net7 vssd1 vssd1 vccd1 vccd1 _0367_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_30_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout119_A net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_59_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_28_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_2_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_15_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_35_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_70_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_42_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_14_Right_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_2_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_78_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_2_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_23_Right_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_78_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_46_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_73_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_92_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_18_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_92_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_32_Right_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_44_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0900_ net102 _0284_ _0288_ _0289_ _0277_ vssd1 vssd1 vccd1 vccd1 _0290_ sky130_fd_sc_hd__o311a_1
XFILLER_41_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0831_ _0211_ _0220_ vssd1 vssd1 vccd1 vccd1 _0221_ sky130_fd_sc_hd__nand2_1
X_0762_ net124 net7 vssd1 vssd1 vccd1 vccd1 _0152_ sky130_fd_sc_hd__and2_1
X_0693_ _0008_ _0009_ _0082_ _0081_ vssd1 vssd1 vccd1 vccd1 _0083_ sky130_fd_sc_hd__o31ai_2
XPHY_EDGE_ROW_41_Right_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_96_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1283__Q clk_divider.rollover_flag vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1314_ clknet_2_2__leaf_clk counter_to_35.next_count\[1\] net122 vssd1 vssd1 vccd1
+ vccd1 count\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_96_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_56_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1245_ _0000_ _0594_ vssd1 vssd1 vccd1 vccd1 _0595_ sky130_fd_sc_hd__or2_1
XFILLER_49_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_64_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1176_ net96 _0534_ _0036_ vssd1 vssd1 vccd1 vccd1 _0535_ sky130_fd_sc_hd__a21o_1
XANTENNA__0854__A net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_50_Right_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_24_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_20_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_15_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_21_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_76_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_101_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_75_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_47_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_101_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_28_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_87_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_15_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_70_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_62_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_41_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_11_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_3_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_3_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_78_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_78_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__0658__B net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1030_ net105 _0415_ vssd1 vssd1 vccd1 vccd1 _0416_ sky130_fd_sc_hd__and2_1
XFILLER_34_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_34_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_61_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0814_ net8 net123 vssd1 vssd1 vccd1 vccd1 _0204_ sky130_fd_sc_hd__xor2_1
Xinput20 prescaler[9] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__buf_1
X_0745_ _0131_ _0132_ vssd1 vssd1 vccd1 vccd1 _0135_ sky130_fd_sc_hd__xor2_1
X_0676_ _0059_ _0065_ vssd1 vssd1 vccd1 vccd1 _0066_ sky130_fd_sc_hd__nand2_1
XFILLER_57_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_96_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1228_ _0578_ _0583_ vssd1 vssd1 vccd1 vccd1 _0584_ sky130_fd_sc_hd__nor2_1
XFILLER_16_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_37_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1159_ clk_divider.count_out\[24\] _0514_ vssd1 vssd1 vccd1 vccd1 _0521_ sky130_fd_sc_hd__nor2_1
XFILLER_80_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout99_A net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_89_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_75_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_18_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1312__RESET_B net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_43_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_31_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_39_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_81_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_66_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_93_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1013_ _0344_ _0401_ vssd1 vssd1 vccd1 vccd1 _0403_ sky130_fd_sc_hd__or2_1
XFILLER_81_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_34_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_62_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_89_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0728_ _0116_ _0117_ vssd1 vssd1 vccd1 vccd1 _0118_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_73_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_4_Right_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0659_ _0005_ _0006_ vssd1 vssd1 vccd1 vccd1 _0049_ sky130_fd_sc_hd__nor2_1
XFILLER_69_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_84_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_57_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_25_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_84_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_53_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_13_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_43_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__0761__B net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_68_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_342 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_48_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_59_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_75_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_84_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_63_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_16_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_16_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_71_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_44_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0671__B net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1195__C1 net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_2_2__f_clk_X clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_35_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_35_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_50_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_13_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_10_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_57_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_79_Right_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_57_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_56_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_26_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_EDGE_ROW_88_Right_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1177__C1 net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_68_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_97_Right_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_36_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0993_ clk_divider.count_out\[11\] _0191_ _0193_ clk_divider.count_out\[10\] _0382_
+ vssd1 vssd1 vccd1 vccd1 _0383_ sky130_fd_sc_hd__o221ai_2
XFILLER_101_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_86_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_67_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_27_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_39_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_27_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_82_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_53_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_50_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_33_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_79_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_TAPCELL_ROW_69_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_65_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_45_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_65_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_61_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_14_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_68_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1261_ _0600_ _0588_ _0022_ net104 vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__and4b_1
XFILLER_49_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xinput7 prescaler[0] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__clkbuf_4
X_1192_ _0191_ clk_divider.next_count\[11\] clk_divider.next_count\[27\] _0299_ vssd1
+ vssd1 vccd1 vccd1 _0550_ sky130_fd_sc_hd__a22o_1
XFILLER_49_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_76_282 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_64_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_64_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_52_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_32_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_9_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_20_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_30_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0976_ _0362_ _0363_ _0364_ _0365_ vssd1 vssd1 vccd1 vccd1 _0366_ sky130_fd_sc_hd__or4bb_1
XFILLER_9_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_101_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_2_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_66_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_35_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_11_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_11_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_7_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_78_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_2_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_78_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_93_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_65_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_19_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_73_252 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_46_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_92_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_33_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_92_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_1_Left_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_61_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0830_ _0218_ _0219_ vssd1 vssd1 vccd1 vccd1 _0220_ sky130_fd_sc_hd__nor2_1
X_0761_ net124 net7 vssd1 vssd1 vccd1 vccd1 _0151_ sky130_fd_sc_hd__nor2_1
X_0692_ _0072_ _0080_ vssd1 vssd1 vccd1 vccd1 _0082_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_47_Left_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1313_ clknet_2_2__leaf_clk counter_to_35.next_count\[0\] net122 vssd1 vssd1 vccd1
+ vccd1 count\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_96_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1244_ net105 count\[1\] net108 _0580_ vssd1 vssd1 vccd1 vccd1 _0594_ sky130_fd_sc_hd__or4_1
XFILLER_56_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1175_ clk_divider.count_out\[27\] _0529_ vssd1 vssd1 vccd1 vccd1 _0534_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_63_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_35_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_56_Left_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_15_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_32_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_21_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0959_ clk_divider.count_out\[19\] _0347_ vssd1 vssd1 vccd1 vccd1 _0349_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_65_Left_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_76_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_87_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_28_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_83_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_74_Left_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_87_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_28_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_15_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_31_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_43_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_83_Left_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_98_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_78_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_78_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_92_Left_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_61_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0813_ _0004_ net19 vssd1 vssd1 vccd1 vccd1 _0203_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_12_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput10 prescaler[12] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__clkbuf_2
X_0744_ _0011_ net124 vssd1 vssd1 vccd1 vccd1 _0134_ sky130_fd_sc_hd__nand2_1
XFILLER_89_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_0675_ _0060_ _0064_ vssd1 vssd1 vccd1 vccd1 _0065_ sky130_fd_sc_hd__xnor2_1
XFILLER_69_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_57_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1227_ count\[4\] _0577_ vssd1 vssd1 vccd1 vccd1 _0583_ sky130_fd_sc_hd__and2_1
XFILLER_65_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1158_ clk_divider.count_out\[24\] _0514_ vssd1 vssd1 vccd1 vccd1 _0520_ sky130_fd_sc_hd__and2_1
XFILLER_80_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1089_ _0458_ _0461_ _0462_ vssd1 vssd1 vccd1 vccd1 _0463_ sky130_fd_sc_hd__a21o_1
XFILLER_20_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_32_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_89_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_16_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_31_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_43_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_8_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_98_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_3_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_94_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_39_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_93_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_47_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1012_ _0344_ _0401_ vssd1 vssd1 vccd1 vccd1 _0402_ sky130_fd_sc_hd__nor2_1
XFILLER_62_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_22_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0727_ _0096_ _0097_ vssd1 vssd1 vccd1 vccd1 _0117_ sky130_fd_sc_hd__xnor2_1
XFILLER_89_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_73_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0658_ _0006_ net17 vssd1 vssd1 vccd1 vccd1 _0048_ sky130_fd_sc_hd__nand2_1
XFILLER_97_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_84_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_27_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_65_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_13_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_25_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_43_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_21_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_23_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_76_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_0_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_59_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_75_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_29_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_16_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_44_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_17_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_16_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_31_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_8_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_3_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_79_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_94_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_47_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_35_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_50_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_62_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_50_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_13_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_50_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_20_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_58_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_57_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_26_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_13_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_41_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_80_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_80_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_44_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0992_ clk_divider.count_out\[9\] _0195_ _0381_ vssd1 vssd1 vccd1 vccd1 _0382_ sky130_fd_sc_hd__o21ba_1
XFILLER_32_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_101_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_27_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_55_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_67_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_42_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_53_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_82_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_81_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_33_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_79_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_92_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_85_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_69_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_45_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_26_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1260_ _0032_ _0581_ _0588_ vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__and3_1
XFILLER_64_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
Xinput8 prescaler[10] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__clkbuf_4
XFILLER_37_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1191_ _0536_ _0539_ _0543_ _0548_ vssd1 vssd1 vccd1 vccd1 _0549_ sky130_fd_sc_hd__or4_1
XFILLER_76_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_49_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_64_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_24_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_64_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_17_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_30_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0975_ clk_divider.count_out\[12\] _0188_ vssd1 vssd1 vccd1 vccd1 _0365_ sky130_fd_sc_hd__nand2_1
XFILLER_10_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_59_206 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_101_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_101_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_2_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_82_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_66_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_38_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_11_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0778__A net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_58_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_46_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_46_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_73_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_46_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_92_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_25_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_41_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_0760_ net17 _0130_ vssd1 vssd1 vccd1 vccd1 _0150_ sky130_fd_sc_hd__xnor2_1
X_0691_ _0072_ _0080_ vssd1 vssd1 vccd1 vccd1 _0081_ sky130_fd_sc_hd__nand2_1
XFILLER_6_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1295__CLK clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_96_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_69_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1312_ clknet_2_2__leaf_clk counter_to_35.next_flag net122 vssd1 vssd1 vccd1 vccd1
+ net21 sky130_fd_sc_hd__dfrtp_1
XFILLER_96_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_84_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1243_ _0022_ _0588_ _0591_ vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__and3_1
XFILLER_2_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_56_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_37_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1174_ clk_divider.count_out\[27\] net92 net90 vssd1 vssd1 vccd1 vccd1 _0533_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_63_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_15_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_43_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout124_A net12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0958_ clk_divider.count_out\[19\] _0347_ vssd1 vssd1 vccd1 vccd1 _0348_ sky130_fd_sc_hd__nand2_1
XFILLER_20_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_21_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0889_ _0277_ _0278_ vssd1 vssd1 vccd1 vccd1 _0279_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_76_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_101_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_68_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_28_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_16_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_87_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_28_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_70_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_30_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_23_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__0812__A2 net18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_11_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_98_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_78_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_38_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_93_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_78_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_66_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_61_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0812_ _0005_ net18 _0064_ _0063_ vssd1 vssd1 vccd1 vccd1 _0202_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_12_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput11 prescaler[13] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__buf_2
XANTENNA__1299__RESET_B net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0743_ _0131_ _0132_ vssd1 vssd1 vccd1 vccd1 _0133_ sky130_fd_sc_hd__nor2_1
X_0674_ _0051_ _0062_ vssd1 vssd1 vccd1 vccd1 _0064_ sky130_fd_sc_hd__xor2_1
XFILLER_88_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_96_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_96_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_69_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1226_ net103 net104 _0581_ vssd1 vssd1 vccd1 vccd1 _0582_ sky130_fd_sc_hd__or3b_1
XFILLER_65_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1157_ clk_divider.count_out\[24\] net92 net90 vssd1 vssd1 vccd1 vccd1 _0519_ sky130_fd_sc_hd__and3_1
XANTENNA__1310__CLK clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1088_ clk_divider.count_out\[12\] net111 net100 vssd1 vssd1 vccd1 vccd1 _0462_ sky130_fd_sc_hd__o21ai_1
XFILLER_80_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_20_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_0_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input1_X net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_48_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_90_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_43_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_7_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_98_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_98_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_3_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_94_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_39_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_93_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_47_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1011_ _0352_ _0355_ _0356_ _0400_ vssd1 vssd1 vccd1 vccd1 _0401_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_17_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_97_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_62_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0726_ _0010_ net13 _0115_ _0113_ vssd1 vssd1 vccd1 vccd1 _0116_ sky130_fd_sc_hd__a31o_1
XFILLER_89_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_73_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0657_ _0007_ net16 _0046_ _0044_ vssd1 vssd1 vccd1 vccd1 _0047_ sky130_fd_sc_hd__a31o_1
XFILLER_97_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_85_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_57_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_72_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1209_ _0330_ clk_divider.next_count\[20\] vssd1 vssd1 vccd1 vccd1 _0567_ sky130_fd_sc_hd__or2_1
XFILLER_25_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_43_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_21_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_23_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_95_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__1234__X _0589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_75_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input17_A prescaler[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_59_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_63_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_16_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_71_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_16_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_17_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_44_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_12_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_33_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_8_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_3_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_100_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_79_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_67_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_12_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_39_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_54_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_50_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_50_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_20_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0709_ _0078_ _0079_ vssd1 vssd1 vccd1 vccd1 _0099_ sky130_fd_sc_hd__xnor2_2
XFILLER_38_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_58_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_58_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input9_A prescaler[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_72_104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_28_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_56_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_13_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_41_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_79_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_49_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_36_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_28_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_32_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0991_ clk_divider.count_out\[10\] _0193_ vssd1 vssd1 vccd1 vccd1 _0381_ sky130_fd_sc_hd__and2_1
XFILLER_74_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_99_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_94_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_27_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_54_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_82_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_53_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_81_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_50_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_33_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_58_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_5_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_69_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_2_3__f_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_76_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1190_ _0544_ _0545_ _0546_ _0547_ vssd1 vssd1 vccd1 vccd1 _0548_ sky130_fd_sc_hd__or4_1
XFILLER_64_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xinput9 prescaler[11] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__clkbuf_2
XFILLER_91_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_36_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_32_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_32_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_30_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0974_ clk_divider.count_out\[13\] _0186_ vssd1 vssd1 vccd1 vccd1 _0364_ sky130_fd_sc_hd__nand2_1
XFILLER_87_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_59_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_2_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_TAPCELL_ROW_66_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_38_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_35_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_35_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_11_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_50_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0778__B net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_18_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_73_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_61_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_92_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_14_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_61_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_14_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_25_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0690_ _0008_ net15 _0079_ _0077_ vssd1 vssd1 vccd1 vccd1 _0080_ sky130_fd_sc_hd__a31o_1
XFILLER_6_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_6_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0688__B net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1311_ clknet_2_0__leaf_clk clk_divider.next_count\[27\] net120 vssd1 vssd1 vccd1
+ vccd1 clk_divider.count_out\[27\] sky130_fd_sc_hd__dfrtp_2
XFILLER_96_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_EDGE_ROW_10_Right_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1242_ _0581_ _0588_ _0591_ vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__and3_1
XFILLER_2_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_2_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1173_ _0528_ _0531_ _0532_ net98 vssd1 vssd1 vccd1 vccd1 clk_divider.next_count\[26\]
+ sky130_fd_sc_hd__o211a_1
XFILLER_92_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_63_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_15_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0957_ _0247_ _0346_ vssd1 vssd1 vccd1 vccd1 _0347_ sky130_fd_sc_hd__xnor2_2
XFILLER_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout117_A net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0888_ _0270_ _0271_ _0276_ vssd1 vssd1 vccd1 vccd1 _0278_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_76_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_46_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_83_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_28_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_87_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_43_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_43_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_62_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_98_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_3_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_93_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_93_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_74_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_36_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput12 prescaler[1] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_12_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0811_ _0003_ _0200_ vssd1 vssd1 vccd1 vccd1 _0201_ sky130_fd_sc_hd__or2_1
X_0742_ net18 _0110_ vssd1 vssd1 vccd1 vccd1 _0132_ sky130_fd_sc_hd__xnor2_1
XFILLER_6_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0673_ _0051_ _0062_ vssd1 vssd1 vccd1 vccd1 _0063_ sky130_fd_sc_hd__nor2_1
XFILLER_42_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_96_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_69_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_84_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1225_ net107 net106 vssd1 vssd1 vccd1 vccd1 _0581_ sky130_fd_sc_hd__and2b_1
XFILLER_37_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_48_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1156_ _0518_ vssd1 vssd1 vccd1 vccd1 clk_divider.next_count\[23\] sky130_fd_sc_hd__inv_2
XFILLER_80_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_65_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_16_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_25_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1087_ net94 _0459_ _0460_ net111 vssd1 vssd1 vccd1 vccd1 _0461_ sky130_fd_sc_hd__o31a_1
XFILLER_40_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_60_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_20_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_4_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_0_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_57_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_28_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_28_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_83_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_56_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1285__CLK clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_7_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_93_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_19_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1010_ _0361_ _0366_ _0399_ vssd1 vssd1 vccd1 vccd1 _0400_ sky130_fd_sc_hd__or3_1
XFILLER_62_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_17_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_22_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_30_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0725_ _0111_ _0112_ vssd1 vssd1 vccd1 vccd1 _0115_ sky130_fd_sc_hd__xor2_1
X_0656_ _0039_ _0043_ vssd1 vssd1 vccd1 vccd1 _0046_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_73_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_97_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_57_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_69_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_84_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1208_ _0011_ clk_divider.next_count\[6\] _0563_ _0564_ _0565_ vssd1 vssd1 vccd1
+ vccd1 _0566_ sky130_fd_sc_hd__a2111o_1
XFILLER_27_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_65_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_38_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_84_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1139_ clk_divider.count_out\[21\] _0498_ vssd1 vssd1 vccd1 vccd1 _0504_ sky130_fd_sc_hd__nor2_1
XFILLER_80_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_40_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_23_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_48_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_59_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_44_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_71_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_31_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_31_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_8_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_8_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_33_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_8_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_89_Left_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__1300__CLK clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__0977__A net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_39_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_94_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_39_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_94_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_47_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_62_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_8_Right_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_22_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_20_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0708_ _0009_ net14 _0097_ _0095_ vssd1 vssd1 vccd1 vccd1 _0098_ sky130_fd_sc_hd__a31o_1
XFILLER_1_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0639_ net108 clk_divider.rollover_flag _0025_ net106 vssd1 vssd1 vccd1 vccd1 _0031_
+ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_39_Right_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__0697__A1 net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_TAPCELL_ROW_28_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_54_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_54_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_41_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_48_Right_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_21_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_79_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_57_Right_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_95_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_0_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_76_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_91_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_66_Right_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_0990_ clk_divider.count_out\[11\] _0191_ vssd1 vssd1 vccd1 vccd1 _0380_ sky130_fd_sc_hd__nand2_1
XFILLER_32_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_44_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_99_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_75_Right_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_39_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_55_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_84_Right_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_47_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_35_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_50_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_33_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_61_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_93_Right_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_92_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_5_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_69_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_58_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_73_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__1241__A _0589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_41_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_101_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_14_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_101_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_39_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_37_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_64_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_91_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_17_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_55_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_44_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_9_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0973_ clk_divider.count_out\[12\] _0188_ vssd1 vssd1 vccd1 vccd1 _0363_ sky130_fd_sc_hd__nor2_1
XFILLER_9_595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_99_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_95_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_2_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_66_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_38_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_70_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_43_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_11_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_51_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_19_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_61_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_14_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1315__RESET_B net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_41_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_69_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_37_6 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1310_ clknet_2_0__leaf_clk clk_divider.next_count\[26\] net120 vssd1 vssd1 vccd1
+ vccd1 clk_divider.count_out\[26\] sky130_fd_sc_hd__dfrtp_1
X_1241_ _0589_ _0593_ vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__nor2_1
XFILLER_1_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_16_Left_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_2_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1172_ clk_divider.count_out\[26\] net110 vssd1 vssd1 vccd1 vccd1 _0532_ sky130_fd_sc_hd__or2_1
XFILLER_92_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_35_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_32_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_25_Left_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0956_ _0242_ _0345_ _0240_ vssd1 vssd1 vccd1 vccd1 _0346_ sky130_fd_sc_hd__a21oi_1
X_0887_ _0270_ _0271_ _0276_ vssd1 vssd1 vccd1 vccd1 _0277_ sky130_fd_sc_hd__nand3_1
XFILLER_101_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_34_Left_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_83_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_28_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_43_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_87_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_24_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_43_Left_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_62_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_7_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_98_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_52_Left_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_59_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_74_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_61_Left_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_30_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
Xinput13 prescaler[2] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_12_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0810_ net11 net125 vssd1 vssd1 vccd1 vccd1 _0200_ sky130_fd_sc_hd__nand2_1
XFILLER_52_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0741_ net17 _0130_ vssd1 vssd1 vccd1 vccd1 _0131_ sky130_fd_sc_hd__nand2_1
X_0672_ net11 _0061_ vssd1 vssd1 vccd1 vccd1 _0062_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_70_Left_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_96_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_96_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_77_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1224_ net107 net1 _0580_ vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__and3_1
XFILLER_92_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_65_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_48_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1155_ _0513_ _0516_ _0517_ vssd1 vssd1 vccd1 vccd1 _0518_ sky130_fd_sc_hd__a21o_1
XFILLER_65_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_25_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_37_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1086_ clk_divider.count_out\[12\] _0455_ vssd1 vssd1 vccd1 vccd1 _0460_ sky130_fd_sc_hd__nor2_1
XFILLER_80_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_52_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_80_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_33_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_32_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_20_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_20_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0939_ _0233_ _0250_ _0253_ vssd1 vssd1 vccd1 vccd1 _0329_ sky130_fd_sc_hd__and3_1
XFILLER_88_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_87_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_57_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_75_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_56_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_71_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
Xclkbuf_2_2__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_2_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_83_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_16_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_43_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_98_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_78_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_93_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_59_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_47_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_47_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_74_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_17_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_45_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_62_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_62_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_15_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_63_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_8_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0724_ _0010_ net13 vssd1 vssd1 vccd1 vccd1 _0114_ sky130_fd_sc_hd__nand2_1
X_0655_ _0007_ net16 vssd1 vssd1 vccd1 vccd1 _0045_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_73_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_97_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_38_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_72_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1207_ _0502_ _0505_ _0506_ _0326_ vssd1 vssd1 vccd1 vccd1 _0565_ sky130_fd_sc_hd__a211oi_1
XFILLER_65_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_53_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_84_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1138_ clk_divider.count_out\[21\] _0498_ vssd1 vssd1 vccd1 vccd1 _0503_ sky130_fd_sc_hd__and2_1
X_1069_ clk_divider.count_out\[9\] _0443_ vssd1 vssd1 vccd1 vccd1 _0446_ sky130_fd_sc_hd__nand2_1
XFILLER_43_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_51_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_95_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_59_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_44_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_56_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_31_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_44_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_8_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_12_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__0977__B net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_67_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_94_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_79_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_54_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_94_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_35_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0707_ _0093_ _0094_ vssd1 vssd1 vccd1 vccd1 _0097_ sky130_fd_sc_hd__xor2_1
XFILLER_89_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_0638_ count\[1\] net108 clk_divider.rollover_flag _0025_ vssd1 vssd1 vccd1 vccd1
+ _0030_ sky130_fd_sc_hd__nand4_1
XFILLER_97_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_85_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_28_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_56_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_13_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__1230__C net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1239__A _0589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_5_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_49_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_36_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_76_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_17_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_8_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_40_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_8_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1298__CLK clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_79_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_39_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_94_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_67_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_53_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_62_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_10_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_33_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_61_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_92_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_98_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_58_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_100_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_69_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_58_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_101_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_101_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_41_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_22_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_1_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_76_220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_39_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_49_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_32_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_32_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_20_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0972_ clk_divider.count_out\[13\] _0186_ vssd1 vssd1 vccd1 vccd1 _0362_ sky130_fd_sc_hd__nor2_1
XFILLER_9_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_TAPCELL_ROW_30_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_78_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1045__C net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_95_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_2_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1313__CLK clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_82_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_35_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_11_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_23_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_2_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_61_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_14_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_25_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_14_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_10_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_6_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_6_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1240_ net103 net106 net107 net104 vssd1 vssd1 vccd1 vccd1 _0593_ sky130_fd_sc_hd__or4bb_1
XFILLER_1_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_77_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1171_ net92 _0529_ _0530_ net109 vssd1 vssd1 vccd1 vccd1 _0531_ sky130_fd_sc_hd__o31ai_1
XTAP_TAPCELL_ROW_63_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_24_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_32_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_60_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_15_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_43_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0955_ _0089_ _0127_ _0175_ _0177_ _0252_ vssd1 vssd1 vccd1 vccd1 _0345_ sky130_fd_sc_hd__a41o_1
XFILLER_9_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0886_ net123 _0275_ _0272_ vssd1 vssd1 vccd1 vccd1 _0276_ sky130_fd_sc_hd__a21bo_1
XFILLER_101_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_87_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_101_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1369_ net116 vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__clkbuf_1
XFILLER_55_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_11_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_98_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_93_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_59_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_74_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_30_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_12_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput14 prescaler[3] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__buf_4
X_0740_ net13 net124 vssd1 vssd1 vccd1 vccd1 _0130_ sky130_fd_sc_hd__xor2_1
X_0671_ net123 net19 vssd1 vssd1 vccd1 vccd1 _0061_ sky130_fd_sc_hd__xor2_1
XFILLER_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_84_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1223_ count\[5\] _0579_ vssd1 vssd1 vccd1 vccd1 _0580_ sky130_fd_sc_hd__nor2_1
XFILLER_28_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_96_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_37_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1154_ clk_divider.count_out\[23\] net109 net98 vssd1 vssd1 vccd1 vccd1 _0517_ sky130_fd_sc_hd__o21ai_1
XFILLER_80_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_25_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1085_ clk_divider.count_out\[12\] clk_divider.count_out\[11\] _0450_ vssd1 vssd1
+ vccd1 vccd1 _0459_ sky130_fd_sc_hd__and3_1
XFILLER_80_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_52_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_33_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA_fanout122_A net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_0938_ _0017_ _0324_ _0325_ vssd1 vssd1 vccd1 vccd1 _0328_ sky130_fd_sc_hd__and3_1
X_0869_ net125 _0004_ _0214_ _0257_ vssd1 vssd1 vccd1 vccd1 _0259_ sky130_fd_sc_hd__o31ai_1
XFILLER_88_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_87_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_28_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_83_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_73_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_28_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_56_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_24_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_7_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_22_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_3_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_17_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_62_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_15_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_30_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_25_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0723_ _0111_ _0112_ vssd1 vssd1 vccd1 vccd1 _0113_ sky130_fd_sc_hd__nor2_1
X_0654_ _0039_ _0043_ vssd1 vssd1 vccd1 vccd1 _0044_ sky130_fd_sc_hd__nor2_1
XFILLER_6_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_84_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1206_ _0189_ _0463_ vssd1 vssd1 vccd1 vccd1 _0564_ sky130_fd_sc_hd__nor2_1
XFILLER_65_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_38_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1137_ clk_divider.count_out\[21\] _0404_ vssd1 vssd1 vccd1 vccd1 _0502_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_84_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_25_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_53_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1068_ clk_divider.count_out\[9\] net94 net91 vssd1 vssd1 vccd1 vccd1 _0445_ sky130_fd_sc_hd__and3_1
XFILLER_33_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_5_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_95_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_0_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_30 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_44_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_44_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_12_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_33_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_22_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_94_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_39_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_58_70 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_94_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_47_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_62_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_35_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_95_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_15_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_30_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0706_ _0009_ net14 vssd1 vssd1 vccd1 vccd1 _0096_ sky130_fd_sc_hd__nand2_1
X_0637_ _0026_ _0029_ vssd1 vssd1 vccd1 vccd1 counter_to_35.next_count\[0\] sky130_fd_sc_hd__nor2_1
XFILLER_97_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_38_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1292__RESET_B net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_38_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_56_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_41_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_80_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_5_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_0_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_76_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_76_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA_input15_A prescaler[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_29_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_91_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_44_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_44_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_8_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_60_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_94_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_10_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_39_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_94_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_23_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_81_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_33_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input7_A prescaler[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_85_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_100_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_69_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_26_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_45_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_81_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_41_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_14_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_5_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_30_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_30_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_76_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_EDGE_ROW_101_Right_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input18_X net18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_91_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0971_ _0357_ _0358_ _0359_ _0360_ vssd1 vssd1 vccd1 vccd1 _0361_ sky130_fd_sc_hd__nand4b_1
XFILLER_71_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_13_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_30_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_99_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_95_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_55_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_82_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_66_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_70_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__0702__A net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_73_202 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1288__CLK clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_41_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_6_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_41_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__0612__A net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_77_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_49_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1170_ clk_divider.count_out\[25\] _0520_ clk_divider.count_out\[26\] vssd1 vssd1
+ vccd1 vccd1 _0530_ sky130_fd_sc_hd__a21oi_1
XFILLER_92_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_77_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_37_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_63_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_20_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_15_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0954_ _0309_ _0313_ _0343_ vssd1 vssd1 vccd1 vccd1 _0344_ sky130_fd_sc_hd__or3_1
X_0885_ _0272_ _0274_ vssd1 vssd1 vccd1 vccd1 _0275_ sky130_fd_sc_hd__and2_1
XFILLER_99_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_101_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1368_ net118 vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__clkbuf_1
XFILLER_95_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_68_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1299_ clknet_2_1__leaf_clk clk_divider.next_count\[15\] net120 vssd1 vssd1 vccd1
+ vccd1 clk_divider.count_out\[15\] sky130_fd_sc_hd__dfrtp_4
XFILLER_55_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_23_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_51_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_11_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_98_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_59_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_19_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_74_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_46_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_19_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_34_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0607__A clk_divider.rollover_flag vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_14_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput15 prescaler[4] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_12_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0670_ _0005_ net18 vssd1 vssd1 vccd1 vccd1 _0060_ sky130_fd_sc_hd__nand2_1
XANTENNA__1303__CLK clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_69_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_2_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1222_ count\[4\] _0577_ vssd1 vssd1 vccd1 vccd1 _0579_ sky130_fd_sc_hd__or2_1
XFILLER_77_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_48_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1153_ net92 _0514_ _0515_ net109 vssd1 vssd1 vccd1 vccd1 _0516_ sky130_fd_sc_hd__o31a_1
XFILLER_92_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_37_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1084_ net97 _0402_ clk_divider.count_out\[12\] vssd1 vssd1 vccd1 vccd1 _0458_ sky130_fd_sc_hd__or3b_1
XFILLER_80_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_33_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_33_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_60_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0937_ _0324_ _0325_ _0017_ vssd1 vssd1 vccd1 vccd1 _0327_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout115_A net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0868_ net125 _0004_ _0214_ _0257_ vssd1 vssd1 vccd1 vccd1 _0258_ sky130_fd_sc_hd__or4_1
X_0799_ _0188_ vssd1 vssd1 vccd1 vccd1 _0189_ sky130_fd_sc_hd__inv_2
XFILLER_0_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_56_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_83_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_71_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_43_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_11_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_51_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_22_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_22_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_3_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_93_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_59_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_74_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_17_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_15_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_15_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_25_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_0722_ net19 _0092_ vssd1 vssd1 vccd1 vccd1 _0112_ sky130_fd_sc_hd__xnor2_1
X_0653_ net9 _0041_ vssd1 vssd1 vccd1 vccd1 _0043_ sky130_fd_sc_hd__xnor2_1
XFILLER_40_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_69_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1205_ _0012_ clk_divider.next_count\[5\] vssd1 vssd1 vccd1 vccd1 _0563_ sky130_fd_sc_hd__and2_1
XFILLER_38_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1136_ _0497_ _0500_ _0501_ net99 vssd1 vssd1 vccd1 vccd1 clk_divider.next_count\[20\]
+ sky130_fd_sc_hd__o211a_1
XFILLER_25_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_53_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_84_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_65_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_25_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_80_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1067_ clk_divider.count_out\[8\] net112 _0441_ _0444_ net100 vssd1 vssd1 vccd1 vccd1
+ clk_divider.next_count\[8\] sky130_fd_sc_hd__o221a_1
XANTENNA__0633__A1 clk_divider.rollover_flag vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_4_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA_fanout118_X net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_76_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_84_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_75_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_44_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_16_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_12_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_12_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_22_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_49_Left_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0620__A net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_58_Left_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_35_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_47_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_62_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_15_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_88_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0705_ _0093_ _0094_ vssd1 vssd1 vccd1 vccd1 _0095_ sky130_fd_sc_hd__nor2_1
X_0636_ net108 clk_divider.rollover_flag _0024_ _0025_ _0027_ vssd1 vssd1 vccd1 vccd1
+ _0029_ sky130_fd_sc_hd__a41o_1
XFILLER_58_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_65_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_53_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1119_ clk_divider.count_out\[18\] _0404_ vssd1 vssd1 vccd1 vccd1 _0487_ sky130_fd_sc_hd__nand2_1
XFILLER_26_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_80_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_17_Right_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_0_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_26_Right_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_95_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_28_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_91_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_76_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_63_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_29_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_27_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_56_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_35_Right_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_60_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_8_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_99_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_4_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_44_Right_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_94_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_67_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_94_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_82_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_35_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_81_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_53_Right_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_33_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_62_Right_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0619_ net124 vssd1 vssd1 vccd1 vccd1 _0012_ sky130_fd_sc_hd__inv_2
XFILLER_100_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_85_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_69_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_26_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_38_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_81_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_71_Right_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_101_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_5_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_80_Right_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_30_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA_fanout98_X net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_39_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_49_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_91_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_17_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_44_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_60_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0970_ clk_divider.count_out\[14\] _0184_ vssd1 vssd1 vccd1 vccd1 _0360_ sky130_fd_sc_hd__or2_1
XFILLER_71_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_30_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_95_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_66_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_38_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_82_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_63_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0702__B net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_46_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_92_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_26_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_42_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_6_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_89_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_49_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_77_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_77_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_37_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_49_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_66_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_92_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_63_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_82_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_15_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_43_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0953_ _0319_ _0320_ _0323_ _0342_ vssd1 vssd1 vccd1 vccd1 _0343_ sky130_fd_sc_hd__or4_1
XFILLER_9_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0884_ _0003_ _0268_ _0273_ vssd1 vssd1 vccd1 vccd1 _0274_ sky130_fd_sc_hd__a21o_1
XFILLER_99_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_68_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1367_ net115 vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__clkbuf_1
XFILLER_95_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_83_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1298_ clknet_2_0__leaf_clk clk_divider.next_count\[14\] net119 vssd1 vssd1 vccd1
+ vccd1 clk_divider.count_out\[14\] sky130_fd_sc_hd__dfrtp_1
XFILLER_24_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_51_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_EDGE_ROW_12_Left_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_98_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_87_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_21_Left_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_86_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_19_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_59_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_100_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_46_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_74_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_15_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_36_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_15_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_14_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_14_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_30_Left_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput16 prescaler[5] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_12_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_6_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1157__C net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_84_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1221_ count\[4\] _0577_ vssd1 vssd1 vccd1 vccd1 _0578_ sky130_fd_sc_hd__nor2_1
XFILLER_77_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_65_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_48_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1152_ clk_divider.count_out\[22\] _0503_ clk_divider.count_out\[23\] vssd1 vssd1
+ vccd1 vccd1 _0515_ sky130_fd_sc_hd__a21oi_1
X_1083_ clk_divider.count_out\[11\] net112 _0454_ _0457_ net100 vssd1 vssd1 vccd1
+ vccd1 clk_divider.next_count\[11\] sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_86_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_33_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_0936_ _0324_ _0325_ vssd1 vssd1 vccd1 vccd1 _0326_ sky130_fd_sc_hd__and2_1
XFILLER_9_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0867_ net11 _0256_ vssd1 vssd1 vccd1 vccd1 _0257_ sky130_fd_sc_hd__xnor2_1
X_0798_ _0172_ _0187_ vssd1 vssd1 vccd1 vccd1 _0188_ sky130_fd_sc_hd__nand2_2
XFILLER_87_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_87_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_68_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_56_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_56_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_71_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_24_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_8_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_11_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_22_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_66_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_47_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1280__Y net80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_47_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__0618__A net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_70_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_63_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_15_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_25_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0721_ net18 _0110_ vssd1 vssd1 vccd1 vccd1 _0111_ sky130_fd_sc_hd__nand2_1
X_0652_ net9 _0041_ vssd1 vssd1 vccd1 vccd1 _0042_ sky130_fd_sc_hd__nand2_1
XFILLER_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_97_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_84_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1204_ _0551_ _0555_ _0559_ _0561_ vssd1 vssd1 vccd1 vccd1 _0562_ sky130_fd_sc_hd__or4_1
XFILLER_38_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1135_ clk_divider.count_out\[20\] net110 vssd1 vssd1 vccd1 vccd1 _0501_ sky130_fd_sc_hd__or2_1
XFILLER_38_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_25_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_80_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1066_ net93 _0442_ _0443_ net112 vssd1 vssd1 vccd1 vccd1 _0444_ sky130_fd_sc_hd__o31ai_1
XFILLER_53_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_33_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_40_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_21_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0919_ clk_divider.count_out\[25\] _0308_ vssd1 vssd1 vccd1 vccd1 _0309_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_95_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_88_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_88_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_29_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_17_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_52_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_12_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_12_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_22_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_72_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_74_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA_output21_A net21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_15_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_22_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_50_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1179__A net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0704_ net20 _0074_ vssd1 vssd1 vccd1 vccd1 _0094_ sky130_fd_sc_hd__xnor2_1
Xmax_cap102 _0265_ vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__buf_1
X_0635_ net118 net5 net3 vssd1 vssd1 vccd1 vccd1 _0028_ sky130_fd_sc_hd__or3b_1
XANTENNA__1316__CLK clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1118_ clk_divider.count_out\[17\] net110 net99 _0486_ vssd1 vssd1 vccd1 vccd1 clk_divider.next_count\[17\]
+ sky130_fd_sc_hd__o211a_1
X_1049_ clk_divider.count_out\[5\] net112 vssd1 vssd1 vccd1 vccd1 _0430_ sky130_fd_sc_hd__or2_1
XFILLER_41_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_53_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_70_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__0721__A net18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_95_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_88_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_28_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_91_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_28_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_44_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_56_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_55_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_44_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_4_Left_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1318__RESET_B net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_99_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_5_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_94_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_94_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_85_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_62_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_35_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_16_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_33_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_92_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0618_ net13 vssd1 vssd1 vccd1 vccd1 _0011_ sky130_fd_sc_hd__inv_2
XFILLER_100_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_100_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_85_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_73_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_26_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_45_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_77_Left_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_81_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_14_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_53_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_81_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_41_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_101_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_5_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_86_Left_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1266__B _0605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_30_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_100_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_89_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA_input20_A prescaler[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_95_Left_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_36_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_91_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_55_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_72_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_60_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_30_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0754__A1 net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1383_ net117 vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__clkbuf_1
XFILLER_27_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_66_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_51_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_50_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_58_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_54_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_26_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_96_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_37_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_92_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_63_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_60_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_82_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_0952_ _0327_ _0328_ _0331_ _0341_ vssd1 vssd1 vccd1 vccd1 _0342_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_15_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_0883_ net11 net9 net8 vssd1 vssd1 vccd1 vccd1 _0273_ sky130_fd_sc_hd__and3b_1
XFILLER_99_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_101_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1366_ net114 vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__clkbuf_1
XFILLER_95_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_68_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1297_ clknet_2_3__leaf_clk clk_divider.next_count\[13\] net122 vssd1 vssd1 vccd1
+ vccd1 clk_divider.count_out\[13\] sky130_fd_sc_hd__dfrtp_1
XFILLER_55_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_36_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_87_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_78_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_19_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_74_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_46_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_36_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_27_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_36_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_42_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_14_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_52_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
Xinput17 prescaler[6] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_12_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_6_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_75_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_96_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1220_ net103 net104 net106 vssd1 vssd1 vccd1 vccd1 _0577_ sky130_fd_sc_hd__or3_1
XFILLER_77_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1151_ clk_divider.count_out\[23\] clk_divider.count_out\[22\] _0503_ vssd1 vssd1
+ vccd1 vccd1 _0514_ sky130_fd_sc_hd__and3_1
XFILLER_92_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_65_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_48_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1082_ net93 _0455_ _0456_ net113 vssd1 vssd1 vccd1 vccd1 _0457_ sky130_fd_sc_hd__o31ai_1
XFILLER_93_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_86_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_60_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0935_ _0231_ _0254_ _0266_ vssd1 vssd1 vccd1 vccd1 _0325_ sky130_fd_sc_hd__or3b_1
XFILLER_9_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0866_ net125 net9 net8 vssd1 vssd1 vccd1 vccd1 _0256_ sky130_fd_sc_hd__o21ba_1
X_0797_ _0163_ _0171_ vssd1 vssd1 vccd1 vccd1 _0187_ sky130_fd_sc_hd__or2_1
XFILLER_87_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_56_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_95_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1380__A net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_71_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_24_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__0636__B1 _0027_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_98_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_22_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__1274__B _0605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_74_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_19_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_74_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_47_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_30_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_42_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_0720_ net14 net13 vssd1 vssd1 vccd1 vccd1 _0110_ sky130_fd_sc_hd__xor2_1
XANTENNA__1168__C net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0651_ net18 net17 vssd1 vssd1 vccd1 vccd1 _0041_ sky130_fd_sc_hd__xor2_1
XFILLER_88_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1203_ _0179_ clk_divider.next_count\[17\] _0507_ _0326_ _0560_ vssd1 vssd1 vccd1
+ vccd1 _0561_ sky130_fd_sc_hd__a221o_1
XFILLER_26_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_38_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1134_ net95 _0498_ _0499_ net110 vssd1 vssd1 vccd1 vccd1 _0500_ sky130_fd_sc_hd__o31ai_1
XFILLER_38_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_53_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1065_ clk_divider.count_out\[8\] clk_divider.count_out\[7\] _0431_ vssd1 vssd1 vccd1
+ vccd1 _0443_ sky130_fd_sc_hd__and3_1
XFILLER_92_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_33_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_fanout120_A net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0918_ _0298_ _0307_ vssd1 vssd1 vccd1 vccd1 _0308_ sky130_fd_sc_hd__nand2_1
X_0849_ net15 _0070_ _0069_ vssd1 vssd1 vccd1 vccd1 _0239_ sky130_fd_sc_hd__a21boi_2
XFILLER_88_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_56_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_29_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_71_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_12_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_8_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1269__B _0605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_35_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_58_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_15_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_30_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_30_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0703_ net19 _0092_ vssd1 vssd1 vccd1 vccd1 _0093_ sky130_fd_sc_hd__nand2_1
XFILLER_7_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_0634_ net5 net3 net1 vssd1 vssd1 vccd1 vccd1 _0027_ sky130_fd_sc_hd__and3b_2
XFILLER_97_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_85_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_38_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_65_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1117_ clk_divider.count_out\[17\] _0404_ _0485_ net96 _0036_ vssd1 vssd1 vccd1 vccd1
+ _0486_ sky130_fd_sc_hd__a221o_1
XFILLER_80_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_53_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1048_ net93 _0427_ _0428_ net112 vssd1 vssd1 vccd1 vccd1 _0429_ sky130_fd_sc_hd__o31ai_1
XFILLER_21_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_EDGE_ROW_3_Right_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1016__B1 _0027_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_0_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_95_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_88_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_0_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_28_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_17_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_71_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_55_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_71_187 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_12_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_44_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_100_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_40_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_5_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_67_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_85_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_82_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0646__X _0036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_31_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_31_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_61_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0617_ net14 vssd1 vssd1 vccd1 vccd1 _0010_ sky130_fd_sc_hd__inv_2
XFILLER_100_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_98_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_69_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1091__C net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_41_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_81_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_41_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_101_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_30_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_89_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_1_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_89_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1173__C1 net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_91_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_64_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input13_A prescaler[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_17_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_32_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_80_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_9_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1306__CLK clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_78_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output81_A net81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1382_ net117 vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__clkbuf_1
XFILLER_96_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_23_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_35_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_50_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_31_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_2_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1383__A net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_76_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_76_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_input5_A la_oenb[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_100_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_100_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_46_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_14_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_41_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_81_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_10_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_89_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_49_257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_92_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_64_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_63_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_17_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_82_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1302__RESET_B net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0951_ clk_divider.count_out\[20\] _0330_ vssd1 vssd1 vccd1 vccd1 _0341_ sky130_fd_sc_hd__nor2_1
XFILLER_60_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_13_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_15_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0882_ _0267_ net11 net8 vssd1 vssd1 vccd1 vccd1 _0272_ sky130_fd_sc_hd__or3b_1
XFILLER_56_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_99_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1365_ net116 vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__clkbuf_1
XFILLER_68_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_95_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_83_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1296_ clknet_2_3__leaf_clk clk_divider.next_count\[12\] net121 vssd1 vssd1 vccd1
+ vccd1 clk_divider.count_out\[12\] sky130_fd_sc_hd__dfrtp_2
XFILLER_23_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_63_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_11_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_3_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_87_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_86_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_74_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_15_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_27_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_36_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_42_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_42_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
Xinput18 prescaler[7] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_12_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_40_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_75_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_97_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_65_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1150_ net96 _0402_ clk_divider.count_out\[23\] vssd1 vssd1 vccd1 vccd1 _0513_ sky130_fd_sc_hd__or3b_1
XFILLER_92_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_77_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_48_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1081_ clk_divider.count_out\[11\] _0450_ vssd1 vssd1 vccd1 vccd1 _0456_ sky130_fd_sc_hd__nor2_1
XFILLER_92_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_93_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_86_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_0934_ _0231_ _0254_ _0266_ vssd1 vssd1 vccd1 vccd1 _0324_ sky130_fd_sc_hd__o21bai_1
XFILLER_9_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_0865_ _0250_ _0253_ _0233_ vssd1 vssd1 vccd1 vccd1 _0255_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_97_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0796_ _0173_ _0185_ vssd1 vssd1 vccd1 vccd1 _0186_ sky130_fd_sc_hd__or2_2
XFILLER_88_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_87_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_68_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_83_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1279_ count\[4\] _0022_ _0032_ _0586_ vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__and4_1
XFILLER_28_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1295__RESET_B net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_24_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_24_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__0724__B net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_7_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0740__A net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_79_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_47_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_59_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_86_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xteam_00_150 vssd1 vssd1 vccd1 vccd1 team_00_150/HI la_data_out[24] sky130_fd_sc_hd__conb_1
XFILLER_19_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_74_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_17_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_25_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0650_ _0006_ _0007_ vssd1 vssd1 vccd1 vccd1 _0040_ sky130_fd_sc_hd__nor2_1
XFILLER_6_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_97_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1202_ _0195_ clk_divider.next_count\[9\] clk_divider.next_count\[26\] _0301_ vssd1
+ vssd1 vccd1 vccd1 _0560_ sky130_fd_sc_hd__o22ai_1
XFILLER_19_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_38_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_92_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1133_ clk_divider.count_out\[19\] _0488_ clk_divider.count_out\[20\] vssd1 vssd1
+ vccd1 vccd1 _0499_ sky130_fd_sc_hd__a21oi_1
XFILLER_65_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1064_ clk_divider.count_out\[7\] _0431_ clk_divider.count_out\[8\] vssd1 vssd1 vccd1
+ vccd1 _0442_ sky130_fd_sc_hd__a21oi_1
XFILLER_53_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_61_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_21_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0917_ net125 _0201_ _0294_ _0296_ vssd1 vssd1 vccd1 vccd1 _0307_ sky130_fd_sc_hd__a211o_1
X_0848_ net16 _0237_ vssd1 vssd1 vccd1 vccd1 _0238_ sky130_fd_sc_hd__xnor2_2
XANTENNA_fanout113_A _0035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0779_ _0167_ _0168_ vssd1 vssd1 vccd1 vccd1 _0169_ sky130_fd_sc_hd__nor2_1
XFILLER_88_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_75_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_29_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_68_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_71_303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_56_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_12_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_EDGE_ROW_18_Left_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_58_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_47_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_35_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_58_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_30_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_90_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0702_ net15 net14 vssd1 vssd1 vccd1 vccd1 _0092_ sky130_fd_sc_hd__xor2_1
XFILLER_99_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0633_ clk_divider.rollover_flag _0025_ net108 vssd1 vssd1 vccd1 vccd1 _0026_ sky130_fd_sc_hd__a21oi_1
XFILLER_97_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_65_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_93_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1116_ _0483_ _0484_ vssd1 vssd1 vccd1 vccd1 _0485_ sky130_fd_sc_hd__nor2_1
XFILLER_80_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1047_ clk_divider.count_out\[4\] _0414_ clk_divider.count_out\[5\] vssd1 vssd1 vccd1
+ vccd1 _0428_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_95_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_76_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_49_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_88_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_29_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_17_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_28_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_27_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_71_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_44_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_12_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_40_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_5_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_4_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_69_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_79_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_7_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_13_Right_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_90_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_22_Right_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_7_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_98_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0616_ net15 vssd1 vssd1 vccd1 vccd1 _0009_ sky130_fd_sc_hd__inv_2
XFILLER_100_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_85_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_31_Right_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_69_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_54_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_41_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_53_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_101_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_40_Right_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_89_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_76_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_76_258 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_76_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_4_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_44_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_80_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_71_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_78_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1381_ net116 vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__clkbuf_1
XFILLER_95_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_66_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_23_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_51_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0690__A2 net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0833__A net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA_clkbuf_0_clk_X clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_100_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_86_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_100_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_86_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_39_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_1_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_26_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_26_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_54_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_10_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_22_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_10_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_1_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_77_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_66_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_60_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_60_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_13_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_20_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0950_ _0306_ _0338_ _0339_ _0303_ vssd1 vssd1 vccd1 vccd1 _0340_ sky130_fd_sc_hd__a211oi_1
XFILLER_60_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_71_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0881_ _0267_ _0268_ _0269_ net8 vssd1 vssd1 vccd1 vccd1 _0271_ sky130_fd_sc_hd__a31o_1
XFILLER_63_5 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_99_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_99_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_68_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_68_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1364_ net114 vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__clkbuf_1
XFILLER_68_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1295_ clknet_2_3__leaf_clk clk_divider.next_count\[11\] net121 vssd1 vssd1 vccd1
+ vccd1 clk_divider.count_out\[11\] sky130_fd_sc_hd__dfrtp_2
XFILLER_83_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_51_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_11_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_78_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_59_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_82_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_15_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_42_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_54_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_27_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_42_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_42_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
Xinput19 prescaler[8] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_12_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_75_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0648__A net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_37_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_92_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_65_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1080_ clk_divider.count_out\[11\] _0450_ vssd1 vssd1 vccd1 vccd1 _0455_ sky130_fd_sc_hd__and2_1
XFILLER_92_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_86_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_33_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0933_ clk_divider.count_out\[22\] _0321_ vssd1 vssd1 vccd1 vccd1 _0323_ sky130_fd_sc_hd__xor2_1
X_0864_ _0250_ _0253_ _0233_ vssd1 vssd1 vccd1 vccd1 _0254_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_97_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0795_ _0148_ _0162_ _0172_ vssd1 vssd1 vccd1 vccd1 _0185_ sky130_fd_sc_hd__and3_1
XFILLER_3_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_95_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1278_ _0032_ _0581_ _0604_ vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__and3_1
XFILLER_83_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_24_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_64_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__0636__A2 clk_divider.rollover_flag vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_24_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_3_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_3_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_93_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_19_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xteam_00_151 vssd1 vssd1 vccd1 vccd1 team_00_151/HI la_data_out[25] sky130_fd_sc_hd__conb_1
Xteam_00_140 vssd1 vssd1 vccd1 vccd1 team_00_140/HI la_data_out[14] sky130_fd_sc_hd__conb_1
XFILLER_74_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_47_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_62_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_34_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_45_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_69_Right_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_8_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__0634__C net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_6_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_78_Right_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1201_ _0556_ _0557_ _0558_ vssd1 vssd1 vccd1 vccd1 _0559_ sky130_fd_sc_hd__or3_1
X_1132_ clk_divider.count_out\[20\] clk_divider.count_out\[19\] _0488_ vssd1 vssd1
+ vccd1 vccd1 _0498_ sky130_fd_sc_hd__and3_1
XFILLER_92_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1063_ clk_divider.count_out\[8\] net93 net90 vssd1 vssd1 vccd1 vccd1 _0441_ sky130_fd_sc_hd__and3_1
XFILLER_65_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_92_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_87_Right_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_61_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1028__C1 net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1043__A2 _0035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0916_ _0302_ _0305_ vssd1 vssd1 vccd1 vccd1 _0306_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_96_Right_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0847_ _0234_ _0235_ vssd1 vssd1 vccd1 vccd1 _0237_ sky130_fd_sc_hd__xor2_2
X_0778_ net15 net7 vssd1 vssd1 vccd1 vccd1 _0168_ sky130_fd_sc_hd__nand2_1
XANTENNA__1291__CLK clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_83_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_71_315 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_16_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_44_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_71_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_17_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_24_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_72_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_90_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_35_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_47_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_74_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_28_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_83_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_30_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_30_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0701_ _0009_ _0010_ vssd1 vssd1 vccd1 vccd1 _0091_ sky130_fd_sc_hd__nor2_1
XFILLER_7_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_94_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0632_ count\[5\] _0021_ vssd1 vssd1 vccd1 vccd1 _0025_ sky130_fd_sc_hd__nand2_1
XFILLER_99_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_97_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_85_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_38_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_57_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_93_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_81_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1115_ clk_divider.count_out\[16\] _0474_ clk_divider.count_out\[17\] vssd1 vssd1
+ vccd1 vccd1 _0484_ sky130_fd_sc_hd__a21oi_1
XFILLER_65_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_53_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1046_ clk_divider.count_out\[5\] clk_divider.count_out\[4\] _0414_ vssd1 vssd1 vccd1
+ vccd1 _0427_ sky130_fd_sc_hd__and3_1
XFILLER_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1016__A2 _0036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_88_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_84_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_17_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_27_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_55_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_71_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_44_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_12_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_40_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_8_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_4_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_4_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_79_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_7_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_75_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_63_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_2_3__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_2_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_90_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_63_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload1_A clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_62_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0615_ net16 vssd1 vssd1 vccd1 vccd1 _0008_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_0_Left_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_37_Left_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_66_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_54_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_38_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1029_ _0030_ _0024_ vssd1 vssd1 vccd1 vccd1 _0415_ sky130_fd_sc_hd__and2b_1
XFILLER_41_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_101_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_46_Left_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_55_Left_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_4_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_17_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_55_21 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_57_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_55_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_80_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_64_Left_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__0987__A1 net12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_91_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_73_Left_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1380_ net118 vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__clkbuf_1
XFILLER_96_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_36_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_82_Left_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_35_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_91_Left_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1289__RESET_B net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_86_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_58_226 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_100_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_100_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_1_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_54_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_37_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_25_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_41_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_10_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_10_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_89_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_1_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_18_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_63_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_32_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_71_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_9_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0880_ net8 _0267_ _0268_ _0269_ vssd1 vssd1 vccd1 vccd1 _0270_ sky130_fd_sc_hd__nand4_2
XFILLER_5_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_99_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_101_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1311__RESET_B net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1363_ net114 vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__clkbuf_1
XFILLER_83_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__0828__B net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1294_ clknet_2_3__leaf_clk clk_divider.next_count\[10\] net121 vssd1 vssd1 vccd1
+ vccd1 clk_divider.count_out\[10\] sky130_fd_sc_hd__dfrtp_1
XFILLER_55_207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_36_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_48_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_23_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_31_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_11_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_86_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_86_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_59_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_46_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_100_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_39_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_42_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_14_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_42_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_12_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_40_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_75_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_65_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_92_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_93_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_18_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_48_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_60_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0932_ _0321_ clk_divider.count_out\[22\] vssd1 vssd1 vccd1 vccd1 _0322_ sky130_fd_sc_hd__nand2b_1
X_0863_ _0240_ _0246_ _0248_ _0252_ _0245_ vssd1 vssd1 vccd1 vccd1 _0253_ sky130_fd_sc_hd__a221oi_2
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0794_ _0147_ _0173_ vssd1 vssd1 vccd1 vccd1 _0184_ sky130_fd_sc_hd__xnor2_2
XFILLER_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__0839__A net18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_3_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_83_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1277_ _0603_ _0604_ vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__and2_1
XFILLER_36_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_12_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_24_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_98_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_3_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA_clkbuf_2_1__f_clk_X clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout120 net121 vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__clkbuf_4
XFILLER_47_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_101_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xteam_00_141 vssd1 vssd1 vccd1 vccd1 team_00_141/HI la_data_out[15] sky130_fd_sc_hd__conb_1
XFILLER_86_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xteam_00_130 vssd1 vssd1 vccd1 vccd1 team_00_130/HI la_data_out[4] sky130_fd_sc_hd__conb_1
Xteam_00_152 vssd1 vssd1 vccd1 vccd1 team_00_152/HI la_data_out[26] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_17_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_42_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_63_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_6_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_97_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_97_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_2_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1200_ _0311_ clk_divider.next_count\[24\] vssd1 vssd1 vccd1 vccd1 _0558_ sky130_fd_sc_hd__and2b_1
XFILLER_77_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_65_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1131_ clk_divider.count_out\[20\] net95 net90 vssd1 vssd1 vccd1 vccd1 _0497_ sky130_fd_sc_hd__and3_1
XFILLER_92_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1062_ _0436_ _0439_ _0440_ net101 vssd1 vssd1 vccd1 vccd1 clk_divider.next_count\[7\]
+ sky130_fd_sc_hd__o211a_1
XFILLER_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_21_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_61_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_99_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0915_ _0014_ _0299_ _0300_ _0303_ _0304_ vssd1 vssd1 vccd1 vccd1 _0305_ sky130_fd_sc_hd__a311o_1
X_0846_ _0234_ _0235_ vssd1 vssd1 vccd1 vccd1 _0236_ sky130_fd_sc_hd__nand2_1
X_0777_ _0153_ _0166_ vssd1 vssd1 vccd1 vccd1 _0167_ sky130_fd_sc_hd__nand2_1
XFILLER_0_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_29_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_68_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_71_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_71_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_24_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_24_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_52_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_22_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_79_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_72_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_79_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_94_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_74_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_47_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_62_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_15_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__0645__C net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_90_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1309__CLK clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0700_ net15 net14 vssd1 vssd1 vccd1 vccd1 _0090_ sky130_fd_sc_hd__nor2_1
X_0631_ _0021_ _0023_ vssd1 vssd1 vccd1 vccd1 _0024_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_94_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_38_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_53_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1114_ clk_divider.count_out\[17\] clk_divider.count_out\[16\] _0474_ vssd1 vssd1
+ vccd1 vccd1 _0483_ sky130_fd_sc_hd__and3_1
XFILLER_93_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_19_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1045_ clk_divider.count_out\[5\] net93 net90 vssd1 vssd1 vccd1 vccd1 _0426_ sky130_fd_sc_hd__and3_1
XFILLER_0_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_34_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_9_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0829_ net123 net19 _0217_ vssd1 vssd1 vccd1 vccd1 _0219_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_27_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_25_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_40_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_4_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_5_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_4_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_79_202 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_4_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_79_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_7_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_35_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_47_132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_75_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_90_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_35_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_90_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_16_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_7_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0614_ net17 vssd1 vssd1 vccd1 vccd1 _0007_ sky130_fd_sc_hd__inv_2
XFILLER_98_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1167__C1 net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_7_Right_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_38_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_26_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_53_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1028_ clk_divider.count_out\[3\] _0412_ _0413_ net98 vssd1 vssd1 vccd1 vccd1 clk_divider.next_count\[3\]
+ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_101_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_22_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_101_Left_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout121_X net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_68_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_29_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_72_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_17_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_80_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_13_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1149__C1 net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_89_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_50_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_31_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_98_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_58_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_100_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_86_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_39_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_73_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_65_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_41_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_54_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_25_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_41_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_10_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_22_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_6_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_66_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_2_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_66_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_18_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA_input11_A prescaler[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_60_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_71_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_43_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_5_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_99_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_95_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1362_ net116 vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__clkbuf_1
XFILLER_68_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_68_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1293_ clknet_2_3__leaf_clk clk_divider.next_count\[9\] net121 vssd1 vssd1 vccd1
+ vccd1 clk_divider.count_out\[9\] sky130_fd_sc_hd__dfrtp_4
XFILLER_83_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_55_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_36_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_48_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_91_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_36_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_23_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_51_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_31_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_11_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_59_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input3_A la_data_in[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_98_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_100_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_86_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_39_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_15_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_42_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_52_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_22_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_89 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_10_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_75_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_77_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_77_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA_input14_X net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_48_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_18_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_33_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0931_ _0283_ _0314_ vssd1 vssd1 vccd1 vccd1 _0321_ sky130_fd_sc_hd__xnor2_2
XFILLER_13_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0862_ _0071_ _0087_ _0251_ vssd1 vssd1 vccd1 vccd1 _0252_ sky130_fd_sc_hd__a21oi_1
X_0793_ _0182_ vssd1 vssd1 vccd1 vccd1 _0183_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_97_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_68_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_68_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1276_ _0602_ _0605_ vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__nor2_1
XFILLER_91_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_22_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_3_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_79_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xfanout121 net122 vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__buf_4
Xfanout110 _0035_ vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__buf_2
XANTENNA_input6_X net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_47_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_101_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xteam_00_131 vssd1 vssd1 vccd1 vccd1 team_00_131/HI la_data_out[5] sky130_fd_sc_hd__conb_1
Xteam_00_142 vssd1 vssd1 vccd1 vccd1 team_00_142/HI la_data_out[16] sky130_fd_sc_hd__conb_1
Xteam_00_153 vssd1 vssd1 vccd1 vccd1 team_00_153/HI la_data_out[27] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_17_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_63_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_70_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_30_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_25_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_12_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_97_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_88_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_88_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1130_ clk_divider.count_out\[19\] net110 _0493_ _0496_ net99 vssd1 vssd1 vccd1 vccd1
+ clk_divider.next_count\[19\] sky130_fd_sc_hd__o221a_1
XFILLER_92_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1061_ clk_divider.count_out\[7\] net113 vssd1 vssd1 vccd1 vccd1 _0440_ sky130_fd_sc_hd__or2_1
XFILLER_92_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_73_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_21_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_33_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_99_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0914_ _0003_ _0297_ _0200_ clk_divider.count_out\[27\] vssd1 vssd1 vccd1 vccd1 _0304_
+ sky130_fd_sc_hd__a211oi_1
X_0845_ _0049_ _0210_ vssd1 vssd1 vccd1 vccd1 _0235_ sky130_fd_sc_hd__xor2_2
X_0776_ _0151_ _0152_ _0008_ vssd1 vssd1 vccd1 vccd1 _0166_ sky130_fd_sc_hd__o21ai_1
XFILLER_88_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_29_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_83_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1259_ _0588_ _0603_ vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__and2_1
XFILLER_37_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_83_188 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_24_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_52_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_22_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_50_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_79_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_58_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_58_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_58_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_54 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_83_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_55_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_43_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_90_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_11_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_7_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_0630_ net106 net107 vssd1 vssd1 vccd1 vccd1 _0023_ sky130_fd_sc_hd__nand2_1
XFILLER_7_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_94_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_66_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_65_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1113_ _0482_ vssd1 vssd1 vccd1 vccd1 clk_divider.next_count\[16\] sky130_fd_sc_hd__inv_2
XFILLER_93_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1044_ _0421_ _0424_ _0425_ vssd1 vssd1 vccd1 vccd1 clk_divider.next_count\[4\] sky130_fd_sc_hd__a21oi_1
XFILLER_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_53_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_34_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_21_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_9_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0828_ net123 net19 _0217_ vssd1 vssd1 vccd1 vccd1 _0218_ sky130_fd_sc_hd__and3_1
X_0759_ _0134_ _0135_ vssd1 vssd1 vccd1 vccd1 _0149_ sky130_fd_sc_hd__xnor2_1
XFILLER_69_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_56_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_84_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_40_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_52_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0762__B net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_40_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_100_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_100_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_40_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_60_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_60_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_4_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_79_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1176__B1 _0036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_69_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_7_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_75_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_63_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_90_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_62_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_50_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1305__RESET_B net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_0613_ net18 vssd1 vssd1 vccd1 vccd1 _0006_ sky130_fd_sc_hd__inv_2
XFILLER_98_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_98_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_98_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_85_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_38_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_93_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_66_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_81_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_34_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1027_ clk_divider.count_out\[0\] clk_divider.count_out\[1\] clk_divider.count_out\[3\]
+ clk_divider.count_out\[2\] vssd1 vssd1 vccd1 vccd1 _0414_ sky130_fd_sc_hd__and4_1
XFILLER_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_22_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_32_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_89_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_1_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_39_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_68_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_57_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_72_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_72_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_13_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_32_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_80_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_9_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_13_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_78_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_91_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_20_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_96_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_95_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_48_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_90_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_35_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_16_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_27_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_65_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_54_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_14_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_25_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_54_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_10_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_9_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_92_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_45_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_82_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_5_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1361_ net115 vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__clkbuf_1
Xoutput80 net80 vssd1 vssd1 vccd1 vccd1 gpio_out[31] sky130_fd_sc_hd__buf_2
X_1292_ clknet_2_1__leaf_clk clk_divider.next_count\[8\] net121 vssd1 vssd1 vccd1
+ vccd1 clk_divider.count_out\[8\] sky130_fd_sc_hd__dfrtp_2
XFILLER_95_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_36_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_76_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_36_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_91_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_62_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_31_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_14_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1294__CLK clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_86_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_100_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_86_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_59_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_86_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_74_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__0639__A2 clk_divider.rollover_flag vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_54_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_52_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_10_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_6_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_75_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_96_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_89_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_77_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_18_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_48_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_18_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_86_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_18_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_20_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0930_ clk_divider.count_out\[23\] _0316_ _0317_ vssd1 vssd1 vccd1 vccd1 _0320_ sky130_fd_sc_hd__and3_1
XFILLER_60_278 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_13_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_0861_ _0071_ _0087_ _0106_ _0107_ vssd1 vssd1 vccd1 vccd1 _0251_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_11_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0792_ _0174_ _0181_ vssd1 vssd1 vccd1 vccd1 _0182_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_97_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_47_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_68_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_EDGE_ROW_79_Left_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_68_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1275_ _0600_ _0604_ _0590_ vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__and3b_1
XFILLER_28_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_56_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_36_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_51_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_88_Left_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout122 net6 vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__buf_4
Xfanout100 net101 vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__buf_2
Xfanout111 net113 vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__buf_2
XFILLER_101_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_47_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_59_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
Xteam_00_132 vssd1 vssd1 vccd1 vccd1 team_00_132/HI la_data_out[6] sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_29_Right_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
Xteam_00_154 vssd1 vssd1 vccd1 vccd1 team_00_154/HI la_data_out[28] sky130_fd_sc_hd__conb_1
Xteam_00_143 vssd1 vssd1 vccd1 vccd1 team_00_143/HI la_data_out[17] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_45_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_42_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_70_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_25_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_38_Right_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_10_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_88_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_97_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_88_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_47_Right_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_80_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1060_ net97 _0437_ _0438_ _0036_ vssd1 vssd1 vccd1 vccd1 _0439_ sky130_fd_sc_hd__a31o_1
XFILLER_92_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_18_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_56_Right_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_99_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0913_ _0200_ _0297_ _0201_ clk_divider.count_out\[27\] vssd1 vssd1 vccd1 vccd1 _0303_
+ sky130_fd_sc_hd__o211a_1
X_0844_ _0040_ _0067_ _0066_ vssd1 vssd1 vccd1 vccd1 _0234_ sky130_fd_sc_hd__a21bo_1
X_0775_ _0155_ _0156_ vssd1 vssd1 vccd1 vccd1 _0165_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_65_Right_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_29_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1258_ net106 net107 net103 net104 vssd1 vssd1 vccd1 vccd1 _0603_ sky130_fd_sc_hd__and4b_1
XFILLER_83_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1189_ _0321_ clk_divider.next_count\[22\] vssd1 vssd1 vccd1 vccd1 _0547_ sky130_fd_sc_hd__xor2_1
XFILLER_24_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_EDGE_ROW_74_Right_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_52_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_22_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_EDGE_ROW_83_Right_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_79_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_72_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_75_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_74_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_TAPCELL_ROW_58_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_74_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_62_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_92_Right_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_83_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_11_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_23_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_7_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_94_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_66_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_2_2__f_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1112_ _0477_ _0480_ _0481_ vssd1 vssd1 vccd1 vccd1 _0482_ sky130_fd_sc_hd__a21o_1
X_1043_ clk_divider.count_out\[4\] _0035_ net99 vssd1 vssd1 vccd1 vccd1 _0425_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_53_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_100_Right_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_34_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0827_ _0212_ _0216_ vssd1 vssd1 vccd1 vccd1 _0217_ sky130_fd_sc_hd__xnor2_1
X_0758_ net7 _0143_ vssd1 vssd1 vccd1 vccd1 _0148_ sky130_fd_sc_hd__xnor2_1
XFILLER_1_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0689_ _0075_ _0076_ vssd1 vssd1 vccd1 vccd1 _0079_ sky130_fd_sc_hd__xor2_2
XFILLER_84_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_69_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_28_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_29_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_56_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_57_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_27_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_100_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_40_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_100_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_60_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_69_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_79_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_69_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_7_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_48_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_35_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_90_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_18_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0612_ net19 vssd1 vssd1 vccd1 vccd1 _0005_ sky130_fd_sc_hd__inv_2
XFILLER_98_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_98_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_100_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_39_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_53_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1026_ clk_divider.count_out\[3\] _0412_ vssd1 vssd1 vccd1 vccd1 _0413_ sky130_fd_sc_hd__nand2_1
XFILLER_22_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_22_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_61_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_32_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_15_Left_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_89_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_69_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_4_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_24_Left_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_68_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_44_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_80_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_13_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_40_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_40_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_33_Left_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_91_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_96_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_95_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_67_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_EDGE_ROW_42_Left_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_48_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_90_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_89_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_90_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_43_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_51_Left_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_98_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_98_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_60_Left_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_37_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_25_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_54_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1009_ _0370_ _0383_ _0398_ _0380_ vssd1 vssd1 vccd1 vccd1 _0399_ sky130_fd_sc_hd__or4b_1
XFILLER_22_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_22_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_41_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_9_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_77_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_17_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_82_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_25_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_15_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_40_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_31_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_5_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1360_ net116 vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__clkbuf_1
Xoutput70 net70 vssd1 vssd1 vccd1 vccd1 gpio_out[22] sky130_fd_sc_hd__buf_2
Xoutput81 net81 vssd1 vssd1 vccd1 vccd1 gpio_out[32] sky130_fd_sc_hd__buf_2
XFILLER_95_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1291_ clknet_2_1__leaf_clk clk_divider.next_count\[7\] net121 vssd1 vssd1 vccd1
+ vccd1 clk_divider.count_out\[7\] sky130_fd_sc_hd__dfrtp_2
XFILLER_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_91_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_62_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_91_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_51_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_51_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_14_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_98_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_100_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_36_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_39_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_54_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_82_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_77_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_2_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_2_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_77_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_77 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_92_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_73_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_18_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_45_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_86_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_33_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_26_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0860_ _0127_ _0175_ _0248_ _0249_ vssd1 vssd1 vccd1 vccd1 _0250_ sky130_fd_sc_hd__nand4_2
XTAP_TAPCELL_ROW_11_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0791_ _0125_ _0126_ vssd1 vssd1 vccd1 vccd1 _0181_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_97_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_95_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_68_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1274_ _0598_ _0605_ vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__nor2_1
XFILLER_83_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_19_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_64_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_91_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_51_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0989_ _0372_ _0378_ _0371_ vssd1 vssd1 vccd1 vccd1 _0379_ sky130_fd_sc_hd__a21o_1
Xfanout101 _0410_ vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__clkbuf_2
Xfanout112 net113 vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__clkbuf_4
XFILLER_59_302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_101_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_86_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
Xfanout123 net20 vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__clkbuf_4
XFILLER_86_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
Xteam_00_133 vssd1 vssd1 vccd1 vccd1 team_00_133/HI la_data_out[7] sky130_fd_sc_hd__conb_1
XFILLER_47_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
Xteam_00_144 vssd1 vssd1 vccd1 vccd1 team_00_144/HI la_data_out[18] sky130_fd_sc_hd__conb_1
Xteam_00_155 vssd1 vssd1 vccd1 vccd1 team_00_155/HI la_data_out[29] sky130_fd_sc_hd__conb_1
XFILLER_27_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_15_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_55_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_70_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_15_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_30_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_7_Left_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_10_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_65_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_77_187 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_65_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_18_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_18_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_46_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_16_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1284__CLK clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_99_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0912_ _0299_ _0300_ _0014_ vssd1 vssd1 vccd1 vccd1 _0302_ sky130_fd_sc_hd__a21oi_1
X_0843_ _0231_ _0232_ vssd1 vssd1 vccd1 vccd1 _0233_ sky130_fd_sc_hd__or2_1
X_0774_ _0152_ _0159_ vssd1 vssd1 vccd1 vccd1 _0164_ sky130_fd_sc_hd__xnor2_1
XFILLER_88_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_68_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1257_ _0589_ _0602_ vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__nor2_1
XFILLER_37_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_83_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1188_ _0308_ clk_divider.next_count\[25\] vssd1 vssd1 vccd1 vccd1 _0546_ sky130_fd_sc_hd__xnor2_1
XFILLER_52_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_22_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_101_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_47_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_47_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_58_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_83_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_55_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_70_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_11_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_30_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_7_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_94_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_97_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_24_6 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_65_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_38_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1111_ clk_divider.count_out\[16\] net109 net98 vssd1 vssd1 vccd1 vccd1 _0481_ sky130_fd_sc_hd__o21ai_1
XFILLER_81_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1042_ net93 _0422_ _0423_ net112 vssd1 vssd1 vccd1 vccd1 _0424_ sky130_fd_sc_hd__o31a_1
XFILLER_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_0_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_61_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_21_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_61_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_21_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0826_ _0213_ _0215_ vssd1 vssd1 vccd1 vccd1 _0216_ sky130_fd_sc_hd__nand2_1
X_0757_ _0144_ _0145_ vssd1 vssd1 vccd1 vccd1 _0147_ sky130_fd_sc_hd__xor2_2
XFILLER_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0688_ _0008_ net15 vssd1 vssd1 vccd1 vccd1 _0078_ sky130_fd_sc_hd__nand2_1
XFILLER_69_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_69_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_84_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_29_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1309_ clknet_2_0__leaf_clk clk_divider.next_count\[25\] net119 vssd1 vssd1 vccd1
+ vccd1 clk_divider.count_out\[25\] sky130_fd_sc_hd__dfrtp_4
XFILLER_84_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_72_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_37_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_44_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_40_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_52_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_40_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_100_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_69_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_79_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_7_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_87_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_85_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_90_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_31_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0611_ net123 vssd1 vssd1 vccd1 vccd1 _0004_ sky130_fd_sc_hd__inv_2
XFILLER_98_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_98_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1314__RESET_B net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_66_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_66_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_81_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1025_ _0412_ net98 _0411_ vssd1 vssd1 vccd1 vccd1 clk_divider.next_count\[2\] sky130_fd_sc_hd__and3b_1
XFILLER_22_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_22_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_61_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_32_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0809_ _0180_ _0182_ _0198_ _0179_ vssd1 vssd1 vccd1 vccd1 _0199_ sky130_fd_sc_hd__and4b_1
XFILLER_89_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_39_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_69_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_29_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_68_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__1231__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_71_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_40_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_71_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_9_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_40_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_78_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_91_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_95_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_29_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_48_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_89_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_90_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_35_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_51_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_90_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_16_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_100_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_6_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_98_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_98_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_66_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_27_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_81_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_81_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1008_ _0371_ _0375_ _0376_ _0397_ vssd1 vssd1 vccd1 vccd1 _0398_ sky130_fd_sc_hd__or4_1
XFILLER_25_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_22_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_34_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_41_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_9_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_77_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_85_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_57_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_17_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_33_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_45_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_40_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_9_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_31_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
Xoutput60 net60 vssd1 vssd1 vccd1 vccd1 gpio_out[13] sky130_fd_sc_hd__buf_2
Xoutput82 net82 vssd1 vssd1 vccd1 vccd1 gpio_out[33] sky130_fd_sc_hd__buf_2
Xoutput71 net71 vssd1 vssd1 vccd1 vccd1 gpio_out[23] sky130_fd_sc_hd__buf_2
X_1290_ clknet_2_1__leaf_clk clk_divider.next_count\[6\] net120 vssd1 vssd1 vccd1
+ vccd1 clk_divider.count_out\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_24_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_91_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_63_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_62_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_16_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_70_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_59_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_67_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_22_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_2_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_77_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_77_89 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_93_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_18_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_86_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_45_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_60_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0790_ _0176_ _0177_ vssd1 vssd1 vccd1 vccd1 _0180_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_11_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_97_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_96_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_95_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1273_ _0597_ _0605_ vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__nor2_1
XFILLER_49_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_83_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_64_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_47_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_24_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_51_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0988_ net13 _0019_ _0374_ _0375_ _0377_ vssd1 vssd1 vccd1 vccd1 _0378_ sky130_fd_sc_hd__o32a_1
XFILLER_99_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
Xfanout113 _0035_ vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_101_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout124 net12 vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__clkbuf_4
XFILLER_59_314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_86_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_74_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input1_A en vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_101_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_86_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
Xteam_00_145 vssd1 vssd1 vccd1 vccd1 team_00_145/HI la_data_out[19] sky130_fd_sc_hd__conb_1
XFILLER_67_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xteam_00_134 vssd1 vssd1 vccd1 vccd1 team_00_134/HI la_data_out[8] sky130_fd_sc_hd__conb_1
Xteam_00_156 vssd1 vssd1 vccd1 vccd1 team_00_156/HI la_data_out[30] sky130_fd_sc_hd__conb_1
XFILLER_55_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_82_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_15_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_27_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_55_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_70_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_23_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_53_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_10_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_6_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_88_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_78_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_2_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_77_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA_input12_X net12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_18_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_46_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_73_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_18_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_37_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_61_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_99_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0911_ _0299_ _0300_ vssd1 vssd1 vccd1 vccd1 _0301_ sky130_fd_sc_hd__nand2_1
X_0842_ _0221_ _0223_ _0230_ vssd1 vssd1 vccd1 vccd1 _0232_ sky130_fd_sc_hd__and3_1
X_0773_ _0160_ _0161_ vssd1 vssd1 vccd1 vccd1 _0163_ sky130_fd_sc_hd__xor2_1
XFILLER_52_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_5_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_96_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_56_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_83_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_17_18 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1256_ _0000_ count\[1\] net108 net105 vssd1 vssd1 vccd1 vccd1 _0602_ sky130_fd_sc_hd__or4b_1
XFILLER_49_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_52_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1187_ _0195_ clk_divider.next_count\[9\] _0463_ _0189_ vssd1 vssd1 vccd1 vccd1 _0545_
+ sky130_fd_sc_hd__a22o_1
XFILLER_37_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_52_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_33_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_52_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_22_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input4_X net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_75_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_101_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_28_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_43_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_15_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_83_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_94_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1110_ net92 _0478_ _0479_ net109 vssd1 vssd1 vccd1 vccd1 _0480_ sky130_fd_sc_hd__o31a_1
XFILLER_93_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_6 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1041_ clk_divider.count_out\[4\] _0414_ vssd1 vssd1 vccd1 vccd1 _0423_ sky130_fd_sc_hd__nor2_1
XFILLER_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_34_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_46_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_21_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_34_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0825_ _0004_ _0214_ vssd1 vssd1 vccd1 vccd1 _0215_ sky130_fd_sc_hd__nand2_1
X_0756_ _0144_ _0145_ vssd1 vssd1 vccd1 vccd1 _0146_ sky130_fd_sc_hd__nor2_1
X_0687_ _0075_ _0076_ vssd1 vssd1 vccd1 vccd1 _0077_ sky130_fd_sc_hd__nor2_1
XFILLER_84_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_29_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_57_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_69_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1308_ clknet_2_0__leaf_clk clk_divider.next_count\[24\] net119 vssd1 vssd1 vccd1
+ vccd1 clk_divider.count_out\[24\] sky130_fd_sc_hd__dfrtp_1
XFILLER_84_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1239_ _0589_ _0592_ vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__nor2_1
XFILLER_25_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_56_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_55_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_87_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_7_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_31_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_7_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0610_ net9 vssd1 vssd1 vccd1 vccd1 _0003_ sky130_fd_sc_hd__inv_2
XFILLER_66_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_39_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_15_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_26_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_66_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_19_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1024_ clk_divider.count_out\[2\] net96 _0408_ vssd1 vssd1 vccd1 vccd1 _0412_ sky130_fd_sc_hd__and3_1
XFILLER_53_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_32_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0808_ _0184_ _0186_ _0197_ vssd1 vssd1 vccd1 vccd1 _0198_ sky130_fd_sc_hd__and3_1
XANTENNA__1297__CLK clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0739_ _0011_ _0012_ vssd1 vssd1 vccd1 vccd1 _0129_ sky130_fd_sc_hd__nor2_1
XFILLER_89_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__0669__A2 net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_57_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_68_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_44_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_13_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_40_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_40_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_91_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_95_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_0_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_88_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_48_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_29_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_89_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_90_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_90_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_43_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_45_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_100_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_80 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_6_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_98_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_6_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_98_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_100_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_86_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_39_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_65_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_81_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1007_ _0012_ clk_divider.count_out\[5\] clk_divider.count_out\[4\] _0013_ _0396_
+ vssd1 vssd1 vccd1 vccd1 _0397_ sky130_fd_sc_hd__a221o_1
XFILLER_22_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_41_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_10_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_41_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_9_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_1_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_89_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_85_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1312__CLK clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_25_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_9_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_40_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_13_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_40_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_99_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput50 net50 vssd1 vssd1 vccd1 vccd1 gpio_oeb[4] sky130_fd_sc_hd__buf_2
Xoutput61 net61 vssd1 vssd1 vccd1 vccd1 gpio_out[14] sky130_fd_sc_hd__buf_2
XFILLER_49_9 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_68_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput83 net83 vssd1 vssd1 vccd1 vccd1 gpio_out[3] sky130_fd_sc_hd__buf_2
Xoutput72 net72 vssd1 vssd1 vccd1 vccd1 gpio_out[24] sky130_fd_sc_hd__buf_2
XFILLER_95_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_63_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_82_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_70_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_59_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_98_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_67_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_82_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_50_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_2_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_2_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_77_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_92_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_9_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_41_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_11_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_39_Left_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_96_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1272_ _0595_ _0605_ vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__nor2_1
XFILLER_95_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_67_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_19_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_48_Left_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_91_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_36_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_20_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0987_ net12 _0020_ _0376_ vssd1 vssd1 vccd1 vccd1 _0377_ sky130_fd_sc_hd__o21a_1
XFILLER_87_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout103 count\[3\] vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__clkbuf_2
XFILLER_99_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
Xfanout114 net117 vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__clkbuf_2
Xfanout125 net10 vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__clkbuf_2
XFILLER_59_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_47_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_101_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_86_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xteam_00_157 vssd1 vssd1 vccd1 vccd1 team_00_157/HI la_data_out[31] sky130_fd_sc_hd__conb_1
Xteam_00_146 vssd1 vssd1 vccd1 vccd1 team_00_146/HI la_data_out[20] sky130_fd_sc_hd__conb_1
Xteam_00_135 vssd1 vssd1 vccd1 vccd1 team_00_135/HI la_data_out[9] sky130_fd_sc_hd__conb_1
XFILLER_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_63_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_70_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_11_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_23_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_53_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_10_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__1291__RESET_B net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_2_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_78_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_77_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_77_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_92_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_16_Right_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_37_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_73_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_18_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_44_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_61_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0910_ net11 _0273_ _0296_ _0268_ vssd1 vssd1 vccd1 vccd1 _0300_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_99_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0841_ _0221_ _0223_ _0230_ vssd1 vssd1 vccd1 vccd1 _0231_ sky130_fd_sc_hd__a21oi_1
X_0772_ _0160_ _0161_ vssd1 vssd1 vccd1 vccd1 _0162_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_25_Right_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_45_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_96_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_69_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1255_ _0600_ _0590_ _0588_ vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__and3b_1
XPHY_EDGE_ROW_34_Right_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1186_ _0180_ _0482_ clk_divider.next_count\[26\] _0301_ vssd1 vssd1 vccd1 vccd1
+ _0544_ sky130_fd_sc_hd__a22o_1
XFILLER_91_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_52_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_52_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_20_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_43_Right_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_58_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_101_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_EDGE_ROW_52_Right_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_70_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_28_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_83_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_43_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_23_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_61_Right_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_70_Right_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_38_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1040_ clk_divider.count_out\[4\] _0414_ vssd1 vssd1 vccd1 vccd1 _0422_ sky130_fd_sc_hd__and2_1
XFILLER_19_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_0_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_73_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0824_ net9 net8 vssd1 vssd1 vccd1 vccd1 _0214_ sky130_fd_sc_hd__nor2_1
X_0755_ net124 _0123_ vssd1 vssd1 vccd1 vccd1 _0145_ sky130_fd_sc_hd__xnor2_2
X_0686_ net8 _0038_ vssd1 vssd1 vccd1 vccd1 _0076_ sky130_fd_sc_hd__xnor2_2
XFILLER_96_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_28_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_29_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1307_ clknet_2_0__leaf_clk clk_divider.next_count\[23\] net119 vssd1 vssd1 vccd1
+ vccd1 clk_divider.count_out\[23\] sky130_fd_sc_hd__dfrtp_1
XFILLER_84_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1238_ net103 net106 net107 net104 vssd1 vssd1 vccd1 vccd1 _0592_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_27_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_55_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1169_ clk_divider.count_out\[26\] clk_divider.count_out\[25\] _0520_ vssd1 vssd1
+ vccd1 vccd1 _0529_ sky130_fd_sc_hd__and3_1
XFILLER_52_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_52_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_7_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_85_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_16_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_62_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_70_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_7_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1021__B1 _0027_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_78_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_38_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_66_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_19_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1023_ net96 _0408_ clk_divider.count_out\[2\] vssd1 vssd1 vccd1 vccd1 _0411_ sky130_fd_sc_hd__a21o_1
XFILLER_53_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_81_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_34_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_46_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_34_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_60_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0807_ _0188_ _0191_ _0193_ _0196_ vssd1 vssd1 vccd1 vccd1 _0197_ sky130_fd_sc_hd__and4_1
XFILLER_89_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0738_ _0122_ _0124_ _0126_ vssd1 vssd1 vccd1 vccd1 _0128_ sky130_fd_sc_hd__a21oi_1
X_0669_ _0006_ net17 _0054_ _0053_ vssd1 vssd1 vccd1 vccd1 _0059_ sky130_fd_sc_hd__a31o_1
XFILLER_39_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_84_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_68_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_2_Right_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_84_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_37_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_13_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_71_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_20_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_91_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_75_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_75_254 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_75_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_48_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_63_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_11_Left_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_89_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_16_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_16_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_31_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_100_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_EDGE_ROW_20_Left_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_98_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_94_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_37_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1006_ clk_divider.count_out\[0\] clk_divider.count_out\[1\] clk_divider.count_out\[3\]
+ clk_divider.count_out\[2\] vssd1 vssd1 vccd1 vccd1 _0396_ sky130_fd_sc_hd__or4_1
XFILLER_22_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_34_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_85_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_85_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_45_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_45_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_60_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_9_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_40_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_5_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xoutput40 net40 vssd1 vssd1 vccd1 vccd1 gpio_oeb[26] sky130_fd_sc_hd__buf_2
Xoutput51 net51 vssd1 vssd1 vccd1 vccd1 gpio_oeb[5] sky130_fd_sc_hd__buf_2
XFILLER_95_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
Xoutput84 net84 vssd1 vssd1 vccd1 vccd1 gpio_out[4] sky130_fd_sc_hd__buf_2
Xoutput73 net73 vssd1 vssd1 vccd1 vccd1 gpio_out[25] sky130_fd_sc_hd__buf_2
Xoutput62 net62 vssd1 vssd1 vccd1 vccd1 gpio_out[15] sky130_fd_sc_hd__buf_2
XFILLER_48_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_76_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1287__CLK clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_70_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_99_Right_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_98_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_86_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_39_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_27_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_82_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_27_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_36_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_42_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_10_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_6_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_77_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_89_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_58_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_85_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_86_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_60_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_41_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_11_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_68_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1271_ _0022_ _0591_ _0604_ vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__and3_1
XFILLER_49_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_49_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_64_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_19_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0986_ clk_divider.count_out\[4\] _0013_ net124 _0020_ vssd1 vssd1 vccd1 vccd1 _0376_
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__1302__CLK clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xfanout104 net105 vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__clkbuf_2
XFILLER_99_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
Xfanout115 net117 vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__buf_1
XFILLER_59_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_47_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
Xteam_00_136 vssd1 vssd1 vccd1 vccd1 team_00_136/HI la_data_out[10] sky130_fd_sc_hd__conb_1
XFILLER_67_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
Xteam_00_147 vssd1 vssd1 vccd1 vccd1 team_00_147/HI la_data_out[21] sky130_fd_sc_hd__conb_1
XFILLER_82_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_63_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_27_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_23_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_42_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_12_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_2_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_5_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_2_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_2_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_93_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_73_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_61_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_33_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_44_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_99_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0840_ net18 _0228_ vssd1 vssd1 vccd1 vccd1 _0230_ sky130_fd_sc_hd__xnor2_1
X_0771_ _0129_ _0139_ vssd1 vssd1 vccd1 vccd1 _0161_ sky130_fd_sc_hd__xnor2_1
XFILLER_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_38_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_96_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_96_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_3_Left_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1254_ _0589_ _0600_ vssd1 vssd1 vccd1 vccd1 _0601_ sky130_fd_sc_hd__or2_1
XFILLER_49_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1185_ clk_divider.next_count\[3\] _0540_ _0541_ _0542_ vssd1 vssd1 vccd1 vccd1 _0543_
+ sky130_fd_sc_hd__or4_1
XFILLER_64_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_91_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_24_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_20_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_20_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0969_ clk_divider.count_out\[14\] _0184_ vssd1 vssd1 vccd1 vccd1 _0359_ sky130_fd_sc_hd__nand2_1
XFILLER_3_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0700__A net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_101_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_75_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_28_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_58_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_43_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_83_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_15_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_70_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_67_Left_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_21_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1265__X _0605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_76_Left_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_78_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_2_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_78_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1144__C net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_138 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_19_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_58_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_73_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_85_Left_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0823_ net8 net123 net9 vssd1 vssd1 vccd1 vccd1 _0213_ sky130_fd_sc_hd__o21ai_1
X_0754_ net7 _0143_ _0142_ vssd1 vssd1 vccd1 vccd1 _0144_ sky130_fd_sc_hd__a21boi_2
XPHY_EDGE_ROW_94_Left_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0685_ net123 _0074_ vssd1 vssd1 vccd1 vccd1 _0075_ sky130_fd_sc_hd__nand2_1
X_1306_ clknet_2_0__leaf_clk clk_divider.next_count\[22\] net119 vssd1 vssd1 vccd1
+ vccd1 clk_divider.count_out\[22\] sky130_fd_sc_hd__dfrtp_2
XFILLER_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1237_ _0000_ net105 vssd1 vssd1 vccd1 vccd1 _0591_ sky130_fd_sc_hd__and2_1
XFILLER_25_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1168_ clk_divider.count_out\[26\] net92 net90 vssd1 vssd1 vccd1 vccd1 _0528_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_55_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_52_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_52_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1099_ clk_divider.count_out\[14\] _0404_ _0470_ net97 _0036_ vssd1 vssd1 vccd1 vccd1
+ _0471_ sky130_fd_sc_hd__a221o_1
XFILLER_60_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_85_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_75_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_18_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_90_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_18_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_70_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_16_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_66_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_93_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1022_ clk_divider.count_out\[1\] _0407_ _0409_ net100 vssd1 vssd1 vccd1 vccd1 clk_divider.next_count\[1\]
+ sky130_fd_sc_hd__o211a_1
XFILLER_19_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_34_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_34_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_61_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_TAPCELL_ROW_32_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0806_ _0011_ _0090_ _0151_ _0195_ vssd1 vssd1 vccd1 vccd1 _0196_ sky130_fd_sc_hd__and4_1
X_0737_ _0125_ _0126_ vssd1 vssd1 vccd1 vccd1 _0127_ sky130_fd_sc_hd__nand2b_1
XFILLER_89_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_0668_ _0007_ _0008_ _0057_ _0056_ vssd1 vssd1 vccd1 vccd1 _0058_ sky130_fd_sc_hd__o31ai_2
XFILLER_97_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_29_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_84_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_68_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_45_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_72_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_25_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_13_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_91_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_0_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_75_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_75_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_63_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_16_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_28_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_16_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_100_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_3_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_79_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_20_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_94_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_39_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_66_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_34_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_50_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_1005_ _0344_ _0393_ _0336_ _0340_ vssd1 vssd1 vccd1 vccd1 _0395_ sky130_fd_sc_hd__o211ai_1
XTAP_TAPCELL_ROW_77_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_45_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_85_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_82_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__1312__Q net21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_40_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_9_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_40_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_21_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput41 net41 vssd1 vssd1 vccd1 vccd1 gpio_oeb[27] sky130_fd_sc_hd__buf_2
Xoutput30 net30 vssd1 vssd1 vccd1 vccd1 gpio_oeb[17] sky130_fd_sc_hd__buf_2
Xoutput52 net52 vssd1 vssd1 vccd1 vccd1 gpio_oeb[6] sky130_fd_sc_hd__buf_2
Xoutput85 net85 vssd1 vssd1 vccd1 vccd1 gpio_out[5] sky130_fd_sc_hd__buf_2
Xoutput63 net63 vssd1 vssd1 vccd1 vccd1 gpio_out[16] sky130_fd_sc_hd__buf_2
Xoutput74 net74 vssd1 vssd1 vccd1 vccd1 gpio_out[26] sky130_fd_sc_hd__buf_2
XFILLER_95_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_0_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_62_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_32_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_71_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_70_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
.ends

